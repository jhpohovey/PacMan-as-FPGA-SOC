/*
    This sprite table was generated using 'conv_to_sv.py'. Find out more here: https://github.com/Atrifex/ECE385-HelperTools
    To use, instantiate this module in your color mapper. The SpriteX input should be connected to
        'ObjectXSize - DistX', where ObjectXSize is the width of your object in pixels along the
        x direction. DistX is the horizontal distance between the DrawX pxiel and the top left corner
        of the object in question, so something like: 'DistX = DrawX - ObjectXPosition' is fine.
        Similarly this goes for SpriteY. Warning: If you don't do this, your image will be flipped along
        the axis you ignored. This is a handy way to flip an image if you need to, though.
 
    In the color mapper, you can then simply do something like:
    module ColorMapper(...)
    ...
    logic [7:0] ObjectR, ObjectG, ObjectB
    parameter ObjectXSize = 10'd10;
    parameter ObjectYSize = 10'd10;
    ...
    always_comb
    ...
         if(ObjectOn == 1'b1)
         begin
             Red = ObjectR
             Green = ObjectG
             Blue = ObjectB
         end
     ...
     ObjectSpriteTable ost(
                           .SpriteX(ObjectXSize - DistX), .SpriteY(ObjectYSize - DistY),
                           .SpriteR(ObjectR), .SpriteG(ObjectG), .SpriteB(ObjectB)
                           );
 
     See the comment at the top of the generation script if you're still confused.
*/
module gameover1(input [9:0] SpriteX, SpriteY,
            output [7:0] SpriteR, SpriteG, SpriteB);

logic [9:0] X_Index, Y_Index;

assign X_Index = SpriteX % 10'd8;
assign Y_Index = SpriteY % 10'd8;
logic [9:0] SpriteTableR;

parameter bit [7:0] SpritePaletteR[4:0] = '{8'd255, 8'd222, 8'd128, 8'd71, 8'd0};

	always_comb
	begin
		SpriteTableR = 10'd0;
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableR = SpriteTableR_0_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableR = SpriteTableR_0_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableR = SpriteTableR_0_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableR = SpriteTableR_0_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableR = SpriteTableR_0_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableR = SpriteTableR_0_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableR = SpriteTableR_0_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableR = SpriteTableR_0_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableR = SpriteTableR_0_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableR = SpriteTableR_0_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableR = SpriteTableR_0_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableR = SpriteTableR_0_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableR = SpriteTableR_0_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_0_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableR = SpriteTableR_0_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableR = SpriteTableR_0_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableR = SpriteTableR_0_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableR = SpriteTableR_0_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableR = SpriteTableR_0_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableR = SpriteTableR_0_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableR = SpriteTableR_0_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableR = SpriteTableR_0_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableR = SpriteTableR_0_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableR = SpriteTableR_0_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableR = SpriteTableR_0_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableR = SpriteTableR_0_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableR = SpriteTableR_0_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableR = SpriteTableR_0_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableR = SpriteTableR_0_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableR = SpriteTableR_0_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableR = SpriteTableR_0_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableR = SpriteTableR_0_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableR = SpriteTableR_0_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableR = SpriteTableR_0_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableR = SpriteTableR_0_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableR = SpriteTableR_0_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableR = SpriteTableR_1_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableR = SpriteTableR_1_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableR = SpriteTableR_1_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableR = SpriteTableR_1_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableR = SpriteTableR_1_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableR = SpriteTableR_1_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableR = SpriteTableR_1_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableR = SpriteTableR_1_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableR = SpriteTableR_1_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableR = SpriteTableR_1_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableR = SpriteTableR_1_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableR = SpriteTableR_1_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableR = SpriteTableR_1_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_1_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableR = SpriteTableR_1_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableR = SpriteTableR_1_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableR = SpriteTableR_1_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableR = SpriteTableR_1_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableR = SpriteTableR_1_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableR = SpriteTableR_1_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableR = SpriteTableR_1_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableR = SpriteTableR_1_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableR = SpriteTableR_1_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableR = SpriteTableR_1_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableR = SpriteTableR_1_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableR = SpriteTableR_1_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableR = SpriteTableR_1_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableR = SpriteTableR_1_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableR = SpriteTableR_1_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableR = SpriteTableR_1_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableR = SpriteTableR_1_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableR = SpriteTableR_1_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableR = SpriteTableR_1_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableR = SpriteTableR_1_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableR = SpriteTableR_1_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableR = SpriteTableR_1_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableR = SpriteTableR_2_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableR = SpriteTableR_2_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableR = SpriteTableR_2_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableR = SpriteTableR_2_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableR = SpriteTableR_2_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableR = SpriteTableR_2_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableR = SpriteTableR_2_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableR = SpriteTableR_2_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableR = SpriteTableR_2_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableR = SpriteTableR_2_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableR = SpriteTableR_2_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableR = SpriteTableR_2_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableR = SpriteTableR_2_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_2_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableR = SpriteTableR_2_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableR = SpriteTableR_2_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableR = SpriteTableR_2_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableR = SpriteTableR_2_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableR = SpriteTableR_2_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableR = SpriteTableR_2_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableR = SpriteTableR_2_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableR = SpriteTableR_2_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableR = SpriteTableR_2_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableR = SpriteTableR_2_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableR = SpriteTableR_2_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableR = SpriteTableR_2_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableR = SpriteTableR_2_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableR = SpriteTableR_2_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableR = SpriteTableR_2_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableR = SpriteTableR_2_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableR = SpriteTableR_2_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableR = SpriteTableR_2_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableR = SpriteTableR_2_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableR = SpriteTableR_2_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableR = SpriteTableR_2_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableR = SpriteTableR_2_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableR = SpriteTableR_3_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableR = SpriteTableR_3_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableR = SpriteTableR_3_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableR = SpriteTableR_3_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableR = SpriteTableR_3_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableR = SpriteTableR_3_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableR = SpriteTableR_3_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableR = SpriteTableR_3_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableR = SpriteTableR_3_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableR = SpriteTableR_3_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableR = SpriteTableR_3_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableR = SpriteTableR_3_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableR = SpriteTableR_3_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_3_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableR = SpriteTableR_3_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableR = SpriteTableR_3_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableR = SpriteTableR_3_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableR = SpriteTableR_3_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableR = SpriteTableR_3_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableR = SpriteTableR_3_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableR = SpriteTableR_3_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableR = SpriteTableR_3_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableR = SpriteTableR_3_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableR = SpriteTableR_3_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableR = SpriteTableR_3_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableR = SpriteTableR_3_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableR = SpriteTableR_3_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableR = SpriteTableR_3_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableR = SpriteTableR_3_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableR = SpriteTableR_3_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableR = SpriteTableR_3_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableR = SpriteTableR_3_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableR = SpriteTableR_3_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableR = SpriteTableR_3_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableR = SpriteTableR_3_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableR = SpriteTableR_3_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableR = SpriteTableR_4_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableR = SpriteTableR_4_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableR = SpriteTableR_4_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableR = SpriteTableR_4_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableR = SpriteTableR_4_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableR = SpriteTableR_4_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableR = SpriteTableR_4_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableR = SpriteTableR_4_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableR = SpriteTableR_4_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableR = SpriteTableR_4_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableR = SpriteTableR_4_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableR = SpriteTableR_4_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableR = SpriteTableR_4_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_4_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableR = SpriteTableR_4_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableR = SpriteTableR_4_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableR = SpriteTableR_4_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableR = SpriteTableR_4_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableR = SpriteTableR_4_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableR = SpriteTableR_4_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableR = SpriteTableR_4_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableR = SpriteTableR_4_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableR = SpriteTableR_4_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableR = SpriteTableR_4_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableR = SpriteTableR_4_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableR = SpriteTableR_4_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableR = SpriteTableR_4_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableR = SpriteTableR_4_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableR = SpriteTableR_4_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableR = SpriteTableR_4_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableR = SpriteTableR_4_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableR = SpriteTableR_4_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableR = SpriteTableR_4_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableR = SpriteTableR_4_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableR = SpriteTableR_4_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableR = SpriteTableR_4_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableR = SpriteTableR_5_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableR = SpriteTableR_5_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableR = SpriteTableR_5_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableR = SpriteTableR_5_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableR = SpriteTableR_5_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableR = SpriteTableR_5_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableR = SpriteTableR_5_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableR = SpriteTableR_5_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableR = SpriteTableR_5_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableR = SpriteTableR_5_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableR = SpriteTableR_5_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableR = SpriteTableR_5_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableR = SpriteTableR_5_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_5_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableR = SpriteTableR_5_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableR = SpriteTableR_5_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableR = SpriteTableR_5_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableR = SpriteTableR_5_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableR = SpriteTableR_5_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableR = SpriteTableR_5_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableR = SpriteTableR_5_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableR = SpriteTableR_5_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableR = SpriteTableR_5_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableR = SpriteTableR_5_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableR = SpriteTableR_5_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableR = SpriteTableR_5_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableR = SpriteTableR_5_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableR = SpriteTableR_5_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableR = SpriteTableR_5_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableR = SpriteTableR_5_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableR = SpriteTableR_5_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableR = SpriteTableR_5_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableR = SpriteTableR_5_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableR = SpriteTableR_5_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableR = SpriteTableR_5_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableR = SpriteTableR_5_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableR = SpriteTableR_6_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableR = SpriteTableR_6_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableR = SpriteTableR_6_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableR = SpriteTableR_6_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableR = SpriteTableR_6_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableR = SpriteTableR_6_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableR = SpriteTableR_6_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableR = SpriteTableR_6_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableR = SpriteTableR_6_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableR = SpriteTableR_6_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableR = SpriteTableR_6_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableR = SpriteTableR_6_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableR = SpriteTableR_6_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_6_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableR = SpriteTableR_6_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableR = SpriteTableR_6_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableR = SpriteTableR_6_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableR = SpriteTableR_6_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableR = SpriteTableR_6_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableR = SpriteTableR_6_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableR = SpriteTableR_6_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableR = SpriteTableR_6_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableR = SpriteTableR_6_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableR = SpriteTableR_6_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableR = SpriteTableR_6_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableR = SpriteTableR_6_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableR = SpriteTableR_6_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableR = SpriteTableR_6_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableR = SpriteTableR_6_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableR = SpriteTableR_6_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableR = SpriteTableR_6_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableR = SpriteTableR_6_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableR = SpriteTableR_6_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableR = SpriteTableR_6_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableR = SpriteTableR_6_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableR = SpriteTableR_6_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableR = SpriteTableR_7_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableR = SpriteTableR_7_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableR = SpriteTableR_7_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableR = SpriteTableR_7_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableR = SpriteTableR_7_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableR = SpriteTableR_7_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableR = SpriteTableR_7_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableR = SpriteTableR_7_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableR = SpriteTableR_7_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableR = SpriteTableR_7_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableR = SpriteTableR_7_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableR = SpriteTableR_7_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableR = SpriteTableR_7_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_7_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableR = SpriteTableR_7_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableR = SpriteTableR_7_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableR = SpriteTableR_7_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableR = SpriteTableR_7_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableR = SpriteTableR_7_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableR = SpriteTableR_7_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableR = SpriteTableR_7_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableR = SpriteTableR_7_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableR = SpriteTableR_7_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableR = SpriteTableR_7_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableR = SpriteTableR_7_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableR = SpriteTableR_7_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableR = SpriteTableR_7_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableR = SpriteTableR_7_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableR = SpriteTableR_7_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableR = SpriteTableR_7_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableR = SpriteTableR_7_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableR = SpriteTableR_7_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableR = SpriteTableR_7_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableR = SpriteTableR_7_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableR = SpriteTableR_7_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableR = SpriteTableR_7_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableR = SpriteTableR_8_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableR = SpriteTableR_8_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableR = SpriteTableR_8_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableR = SpriteTableR_8_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableR = SpriteTableR_8_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableR = SpriteTableR_8_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableR = SpriteTableR_8_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableR = SpriteTableR_8_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableR = SpriteTableR_8_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableR = SpriteTableR_8_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableR = SpriteTableR_8_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableR = SpriteTableR_8_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableR = SpriteTableR_8_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_8_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableR = SpriteTableR_8_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableR = SpriteTableR_8_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableR = SpriteTableR_8_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableR = SpriteTableR_8_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableR = SpriteTableR_8_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableR = SpriteTableR_8_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableR = SpriteTableR_8_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableR = SpriteTableR_8_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableR = SpriteTableR_8_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableR = SpriteTableR_8_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableR = SpriteTableR_8_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableR = SpriteTableR_8_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableR = SpriteTableR_8_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableR = SpriteTableR_8_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableR = SpriteTableR_8_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableR = SpriteTableR_8_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableR = SpriteTableR_8_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableR = SpriteTableR_8_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableR = SpriteTableR_8_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableR = SpriteTableR_8_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableR = SpriteTableR_8_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableR = SpriteTableR_8_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableR = SpriteTableR_9_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableR = SpriteTableR_9_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableR = SpriteTableR_9_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableR = SpriteTableR_9_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableR = SpriteTableR_9_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableR = SpriteTableR_9_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableR = SpriteTableR_9_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableR = SpriteTableR_9_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableR = SpriteTableR_9_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableR = SpriteTableR_9_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableR = SpriteTableR_9_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableR = SpriteTableR_9_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableR = SpriteTableR_9_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_9_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableR = SpriteTableR_9_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableR = SpriteTableR_9_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableR = SpriteTableR_9_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableR = SpriteTableR_9_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableR = SpriteTableR_9_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableR = SpriteTableR_9_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableR = SpriteTableR_9_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableR = SpriteTableR_9_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableR = SpriteTableR_9_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableR = SpriteTableR_9_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableR = SpriteTableR_9_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableR = SpriteTableR_9_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableR = SpriteTableR_9_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableR = SpriteTableR_9_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableR = SpriteTableR_9_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableR = SpriteTableR_9_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableR = SpriteTableR_9_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableR = SpriteTableR_9_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableR = SpriteTableR_9_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableR = SpriteTableR_9_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableR = SpriteTableR_9_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableR = SpriteTableR_9_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableR = SpriteTableR_10_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableR = SpriteTableR_10_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableR = SpriteTableR_10_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableR = SpriteTableR_10_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableR = SpriteTableR_10_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableR = SpriteTableR_10_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableR = SpriteTableR_10_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableR = SpriteTableR_10_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableR = SpriteTableR_10_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableR = SpriteTableR_10_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableR = SpriteTableR_10_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableR = SpriteTableR_10_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableR = SpriteTableR_10_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_10_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableR = SpriteTableR_10_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableR = SpriteTableR_10_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableR = SpriteTableR_10_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableR = SpriteTableR_10_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableR = SpriteTableR_10_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableR = SpriteTableR_10_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableR = SpriteTableR_10_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableR = SpriteTableR_10_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableR = SpriteTableR_10_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableR = SpriteTableR_10_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableR = SpriteTableR_10_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableR = SpriteTableR_10_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableR = SpriteTableR_10_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableR = SpriteTableR_10_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableR = SpriteTableR_10_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableR = SpriteTableR_10_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableR = SpriteTableR_10_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableR = SpriteTableR_10_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableR = SpriteTableR_10_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableR = SpriteTableR_10_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableR = SpriteTableR_10_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableR = SpriteTableR_10_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableR = SpriteTableR_11_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableR = SpriteTableR_11_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableR = SpriteTableR_11_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableR = SpriteTableR_11_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableR = SpriteTableR_11_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableR = SpriteTableR_11_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableR = SpriteTableR_11_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableR = SpriteTableR_11_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableR = SpriteTableR_11_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableR = SpriteTableR_11_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableR = SpriteTableR_11_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableR = SpriteTableR_11_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableR = SpriteTableR_11_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_11_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableR = SpriteTableR_11_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableR = SpriteTableR_11_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableR = SpriteTableR_11_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableR = SpriteTableR_11_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableR = SpriteTableR_11_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableR = SpriteTableR_11_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableR = SpriteTableR_11_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableR = SpriteTableR_11_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableR = SpriteTableR_11_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableR = SpriteTableR_11_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableR = SpriteTableR_11_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableR = SpriteTableR_11_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableR = SpriteTableR_11_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableR = SpriteTableR_11_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableR = SpriteTableR_11_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableR = SpriteTableR_11_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableR = SpriteTableR_11_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableR = SpriteTableR_11_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableR = SpriteTableR_11_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableR = SpriteTableR_11_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableR = SpriteTableR_11_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableR = SpriteTableR_11_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableR = SpriteTableR_12_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableR = SpriteTableR_12_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableR = SpriteTableR_12_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableR = SpriteTableR_12_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableR = SpriteTableR_12_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableR = SpriteTableR_12_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableR = SpriteTableR_12_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableR = SpriteTableR_12_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableR = SpriteTableR_12_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableR = SpriteTableR_12_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableR = SpriteTableR_12_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableR = SpriteTableR_12_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableR = SpriteTableR_12_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_12_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableR = SpriteTableR_12_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableR = SpriteTableR_12_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableR = SpriteTableR_12_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableR = SpriteTableR_12_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableR = SpriteTableR_12_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableR = SpriteTableR_12_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableR = SpriteTableR_12_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableR = SpriteTableR_12_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableR = SpriteTableR_12_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableR = SpriteTableR_12_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableR = SpriteTableR_12_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableR = SpriteTableR_12_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableR = SpriteTableR_12_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableR = SpriteTableR_12_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableR = SpriteTableR_12_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableR = SpriteTableR_12_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableR = SpriteTableR_12_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableR = SpriteTableR_12_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableR = SpriteTableR_12_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableR = SpriteTableR_12_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableR = SpriteTableR_12_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableR = SpriteTableR_12_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableR = SpriteTableR_13_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableR = SpriteTableR_13_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableR = SpriteTableR_13_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableR = SpriteTableR_13_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableR = SpriteTableR_13_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableR = SpriteTableR_13_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableR = SpriteTableR_13_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableR = SpriteTableR_13_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableR = SpriteTableR_13_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableR = SpriteTableR_13_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableR = SpriteTableR_13_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableR = SpriteTableR_13_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableR = SpriteTableR_13_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_13_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableR = SpriteTableR_13_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableR = SpriteTableR_13_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableR = SpriteTableR_13_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableR = SpriteTableR_13_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableR = SpriteTableR_13_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableR = SpriteTableR_13_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableR = SpriteTableR_13_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableR = SpriteTableR_13_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableR = SpriteTableR_13_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableR = SpriteTableR_13_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableR = SpriteTableR_13_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableR = SpriteTableR_13_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableR = SpriteTableR_13_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableR = SpriteTableR_13_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableR = SpriteTableR_13_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableR = SpriteTableR_13_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableR = SpriteTableR_13_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableR = SpriteTableR_13_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableR = SpriteTableR_13_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableR = SpriteTableR_13_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableR = SpriteTableR_13_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableR = SpriteTableR_13_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableR = SpriteTableR_14_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableR = SpriteTableR_14_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableR = SpriteTableR_14_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableR = SpriteTableR_14_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableR = SpriteTableR_14_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableR = SpriteTableR_14_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableR = SpriteTableR_14_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableR = SpriteTableR_14_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableR = SpriteTableR_14_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableR = SpriteTableR_14_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableR = SpriteTableR_14_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableR = SpriteTableR_14_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableR = SpriteTableR_14_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_14_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableR = SpriteTableR_14_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableR = SpriteTableR_14_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableR = SpriteTableR_14_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableR = SpriteTableR_14_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableR = SpriteTableR_14_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableR = SpriteTableR_14_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableR = SpriteTableR_14_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableR = SpriteTableR_14_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableR = SpriteTableR_14_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableR = SpriteTableR_14_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableR = SpriteTableR_14_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableR = SpriteTableR_14_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableR = SpriteTableR_14_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableR = SpriteTableR_14_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableR = SpriteTableR_14_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableR = SpriteTableR_14_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableR = SpriteTableR_14_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableR = SpriteTableR_14_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableR = SpriteTableR_14_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableR = SpriteTableR_14_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableR = SpriteTableR_14_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableR = SpriteTableR_14_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableR = SpriteTableR_15_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableR = SpriteTableR_15_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableR = SpriteTableR_15_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableR = SpriteTableR_15_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableR = SpriteTableR_15_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableR = SpriteTableR_15_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableR = SpriteTableR_15_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableR = SpriteTableR_15_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableR = SpriteTableR_15_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableR = SpriteTableR_15_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableR = SpriteTableR_15_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableR = SpriteTableR_15_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableR = SpriteTableR_15_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_15_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableR = SpriteTableR_15_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableR = SpriteTableR_15_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableR = SpriteTableR_15_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableR = SpriteTableR_15_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableR = SpriteTableR_15_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableR = SpriteTableR_15_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableR = SpriteTableR_15_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableR = SpriteTableR_15_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableR = SpriteTableR_15_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableR = SpriteTableR_15_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableR = SpriteTableR_15_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableR = SpriteTableR_15_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableR = SpriteTableR_15_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableR = SpriteTableR_15_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableR = SpriteTableR_15_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableR = SpriteTableR_15_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableR = SpriteTableR_15_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableR = SpriteTableR_15_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableR = SpriteTableR_15_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableR = SpriteTableR_15_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableR = SpriteTableR_15_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableR = SpriteTableR_15_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableR = SpriteTableR_16_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableR = SpriteTableR_16_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableR = SpriteTableR_16_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableR = SpriteTableR_16_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableR = SpriteTableR_16_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableR = SpriteTableR_16_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableR = SpriteTableR_16_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableR = SpriteTableR_16_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableR = SpriteTableR_16_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableR = SpriteTableR_16_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableR = SpriteTableR_16_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableR = SpriteTableR_16_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableR = SpriteTableR_16_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_16_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableR = SpriteTableR_16_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableR = SpriteTableR_16_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableR = SpriteTableR_16_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableR = SpriteTableR_16_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableR = SpriteTableR_16_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableR = SpriteTableR_16_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableR = SpriteTableR_16_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableR = SpriteTableR_16_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableR = SpriteTableR_16_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableR = SpriteTableR_16_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableR = SpriteTableR_16_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableR = SpriteTableR_16_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableR = SpriteTableR_16_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableR = SpriteTableR_16_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableR = SpriteTableR_16_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableR = SpriteTableR_16_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableR = SpriteTableR_16_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableR = SpriteTableR_16_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableR = SpriteTableR_16_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableR = SpriteTableR_16_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableR = SpriteTableR_16_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableR = SpriteTableR_16_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableR = SpriteTableR_17_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableR = SpriteTableR_17_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableR = SpriteTableR_17_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableR = SpriteTableR_17_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableR = SpriteTableR_17_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableR = SpriteTableR_17_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableR = SpriteTableR_17_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableR = SpriteTableR_17_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableR = SpriteTableR_17_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableR = SpriteTableR_17_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableR = SpriteTableR_17_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableR = SpriteTableR_17_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableR = SpriteTableR_17_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_17_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableR = SpriteTableR_17_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableR = SpriteTableR_17_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableR = SpriteTableR_17_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableR = SpriteTableR_17_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableR = SpriteTableR_17_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableR = SpriteTableR_17_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableR = SpriteTableR_17_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableR = SpriteTableR_17_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableR = SpriteTableR_17_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableR = SpriteTableR_17_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableR = SpriteTableR_17_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableR = SpriteTableR_17_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableR = SpriteTableR_17_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableR = SpriteTableR_17_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableR = SpriteTableR_17_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableR = SpriteTableR_17_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableR = SpriteTableR_17_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableR = SpriteTableR_17_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableR = SpriteTableR_17_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableR = SpriteTableR_17_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableR = SpriteTableR_17_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableR = SpriteTableR_17_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableR = SpriteTableR_18_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableR = SpriteTableR_18_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableR = SpriteTableR_18_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableR = SpriteTableR_18_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableR = SpriteTableR_18_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableR = SpriteTableR_18_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableR = SpriteTableR_18_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableR = SpriteTableR_18_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableR = SpriteTableR_18_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableR = SpriteTableR_18_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableR = SpriteTableR_18_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableR = SpriteTableR_18_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableR = SpriteTableR_18_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_18_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableR = SpriteTableR_18_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableR = SpriteTableR_18_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableR = SpriteTableR_18_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableR = SpriteTableR_18_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableR = SpriteTableR_18_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableR = SpriteTableR_18_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableR = SpriteTableR_18_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableR = SpriteTableR_18_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableR = SpriteTableR_18_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableR = SpriteTableR_18_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableR = SpriteTableR_18_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableR = SpriteTableR_18_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableR = SpriteTableR_18_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableR = SpriteTableR_18_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableR = SpriteTableR_18_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableR = SpriteTableR_18_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableR = SpriteTableR_18_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableR = SpriteTableR_18_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableR = SpriteTableR_18_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableR = SpriteTableR_18_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableR = SpriteTableR_18_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableR = SpriteTableR_18_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableR = SpriteTableR_19_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableR = SpriteTableR_19_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableR = SpriteTableR_19_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableR = SpriteTableR_19_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableR = SpriteTableR_19_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableR = SpriteTableR_19_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableR = SpriteTableR_19_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableR = SpriteTableR_19_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableR = SpriteTableR_19_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableR = SpriteTableR_19_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableR = SpriteTableR_19_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableR = SpriteTableR_19_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableR = SpriteTableR_19_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_19_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableR = SpriteTableR_19_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableR = SpriteTableR_19_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableR = SpriteTableR_19_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableR = SpriteTableR_19_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableR = SpriteTableR_19_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableR = SpriteTableR_19_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableR = SpriteTableR_19_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableR = SpriteTableR_19_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableR = SpriteTableR_19_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableR = SpriteTableR_19_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableR = SpriteTableR_19_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableR = SpriteTableR_19_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableR = SpriteTableR_19_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableR = SpriteTableR_19_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableR = SpriteTableR_19_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableR = SpriteTableR_19_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableR = SpriteTableR_19_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableR = SpriteTableR_19_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableR = SpriteTableR_19_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableR = SpriteTableR_19_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableR = SpriteTableR_19_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableR = SpriteTableR_19_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableR = SpriteTableR_20_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableR = SpriteTableR_20_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableR = SpriteTableR_20_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableR = SpriteTableR_20_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableR = SpriteTableR_20_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableR = SpriteTableR_20_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableR = SpriteTableR_20_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableR = SpriteTableR_20_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableR = SpriteTableR_20_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableR = SpriteTableR_20_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableR = SpriteTableR_20_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableR = SpriteTableR_20_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableR = SpriteTableR_20_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_20_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableR = SpriteTableR_20_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableR = SpriteTableR_20_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableR = SpriteTableR_20_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableR = SpriteTableR_20_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableR = SpriteTableR_20_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableR = SpriteTableR_20_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableR = SpriteTableR_20_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableR = SpriteTableR_20_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableR = SpriteTableR_20_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableR = SpriteTableR_20_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableR = SpriteTableR_20_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableR = SpriteTableR_20_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableR = SpriteTableR_20_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableR = SpriteTableR_20_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableR = SpriteTableR_20_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableR = SpriteTableR_20_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableR = SpriteTableR_20_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableR = SpriteTableR_20_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableR = SpriteTableR_20_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableR = SpriteTableR_20_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableR = SpriteTableR_20_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableR = SpriteTableR_20_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableR = SpriteTableR_21_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableR = SpriteTableR_21_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableR = SpriteTableR_21_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableR = SpriteTableR_21_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableR = SpriteTableR_21_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableR = SpriteTableR_21_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableR = SpriteTableR_21_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableR = SpriteTableR_21_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableR = SpriteTableR_21_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableR = SpriteTableR_21_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableR = SpriteTableR_21_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableR = SpriteTableR_21_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableR = SpriteTableR_21_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_21_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableR = SpriteTableR_21_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableR = SpriteTableR_21_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableR = SpriteTableR_21_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableR = SpriteTableR_21_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableR = SpriteTableR_21_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableR = SpriteTableR_21_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableR = SpriteTableR_21_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableR = SpriteTableR_21_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableR = SpriteTableR_21_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableR = SpriteTableR_21_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableR = SpriteTableR_21_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableR = SpriteTableR_21_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableR = SpriteTableR_21_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableR = SpriteTableR_21_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableR = SpriteTableR_21_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableR = SpriteTableR_21_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableR = SpriteTableR_21_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableR = SpriteTableR_21_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableR = SpriteTableR_21_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableR = SpriteTableR_21_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableR = SpriteTableR_21_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableR = SpriteTableR_21_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableR = SpriteTableR_22_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableR = SpriteTableR_22_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableR = SpriteTableR_22_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableR = SpriteTableR_22_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableR = SpriteTableR_22_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableR = SpriteTableR_22_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableR = SpriteTableR_22_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableR = SpriteTableR_22_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableR = SpriteTableR_22_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableR = SpriteTableR_22_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableR = SpriteTableR_22_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableR = SpriteTableR_22_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableR = SpriteTableR_22_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_22_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableR = SpriteTableR_22_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableR = SpriteTableR_22_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableR = SpriteTableR_22_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableR = SpriteTableR_22_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableR = SpriteTableR_22_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableR = SpriteTableR_22_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableR = SpriteTableR_22_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableR = SpriteTableR_22_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableR = SpriteTableR_22_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableR = SpriteTableR_22_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableR = SpriteTableR_22_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableR = SpriteTableR_22_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableR = SpriteTableR_22_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableR = SpriteTableR_22_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableR = SpriteTableR_22_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableR = SpriteTableR_22_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableR = SpriteTableR_22_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableR = SpriteTableR_22_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableR = SpriteTableR_22_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableR = SpriteTableR_22_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableR = SpriteTableR_22_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableR = SpriteTableR_22_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableR = SpriteTableR_23_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableR = SpriteTableR_23_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableR = SpriteTableR_23_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableR = SpriteTableR_23_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableR = SpriteTableR_23_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableR = SpriteTableR_23_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableR = SpriteTableR_23_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableR = SpriteTableR_23_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableR = SpriteTableR_23_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableR = SpriteTableR_23_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableR = SpriteTableR_23_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableR = SpriteTableR_23_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableR = SpriteTableR_23_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_23_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableR = SpriteTableR_23_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableR = SpriteTableR_23_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableR = SpriteTableR_23_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableR = SpriteTableR_23_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableR = SpriteTableR_23_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableR = SpriteTableR_23_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableR = SpriteTableR_23_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableR = SpriteTableR_23_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableR = SpriteTableR_23_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableR = SpriteTableR_23_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableR = SpriteTableR_23_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableR = SpriteTableR_23_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableR = SpriteTableR_23_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableR = SpriteTableR_23_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableR = SpriteTableR_23_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableR = SpriteTableR_23_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableR = SpriteTableR_23_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableR = SpriteTableR_23_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableR = SpriteTableR_23_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableR = SpriteTableR_23_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableR = SpriteTableR_23_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableR = SpriteTableR_23_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableR = SpriteTableR_24_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableR = SpriteTableR_24_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableR = SpriteTableR_24_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableR = SpriteTableR_24_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableR = SpriteTableR_24_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableR = SpriteTableR_24_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableR = SpriteTableR_24_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableR = SpriteTableR_24_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableR = SpriteTableR_24_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableR = SpriteTableR_24_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableR = SpriteTableR_24_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableR = SpriteTableR_24_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableR = SpriteTableR_24_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_24_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableR = SpriteTableR_24_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableR = SpriteTableR_24_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableR = SpriteTableR_24_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableR = SpriteTableR_24_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableR = SpriteTableR_24_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableR = SpriteTableR_24_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableR = SpriteTableR_24_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableR = SpriteTableR_24_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableR = SpriteTableR_24_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableR = SpriteTableR_24_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableR = SpriteTableR_24_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableR = SpriteTableR_24_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableR = SpriteTableR_24_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableR = SpriteTableR_24_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableR = SpriteTableR_24_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableR = SpriteTableR_24_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableR = SpriteTableR_24_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableR = SpriteTableR_24_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableR = SpriteTableR_24_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableR = SpriteTableR_24_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableR = SpriteTableR_24_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableR = SpriteTableR_24_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableR = SpriteTableR_25_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableR = SpriteTableR_25_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableR = SpriteTableR_25_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableR = SpriteTableR_25_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableR = SpriteTableR_25_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableR = SpriteTableR_25_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableR = SpriteTableR_25_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableR = SpriteTableR_25_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableR = SpriteTableR_25_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableR = SpriteTableR_25_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableR = SpriteTableR_25_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableR = SpriteTableR_25_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableR = SpriteTableR_25_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_25_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableR = SpriteTableR_25_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableR = SpriteTableR_25_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableR = SpriteTableR_25_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableR = SpriteTableR_25_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableR = SpriteTableR_25_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableR = SpriteTableR_25_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableR = SpriteTableR_25_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableR = SpriteTableR_25_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableR = SpriteTableR_25_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableR = SpriteTableR_25_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableR = SpriteTableR_25_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableR = SpriteTableR_25_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableR = SpriteTableR_25_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableR = SpriteTableR_25_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableR = SpriteTableR_25_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableR = SpriteTableR_25_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableR = SpriteTableR_25_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableR = SpriteTableR_25_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableR = SpriteTableR_25_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableR = SpriteTableR_25_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableR = SpriteTableR_25_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableR = SpriteTableR_25_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableR = SpriteTableR_26_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableR = SpriteTableR_26_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableR = SpriteTableR_26_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableR = SpriteTableR_26_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableR = SpriteTableR_26_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableR = SpriteTableR_26_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableR = SpriteTableR_26_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableR = SpriteTableR_26_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableR = SpriteTableR_26_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableR = SpriteTableR_26_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableR = SpriteTableR_26_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableR = SpriteTableR_26_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableR = SpriteTableR_26_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_26_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableR = SpriteTableR_26_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableR = SpriteTableR_26_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableR = SpriteTableR_26_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableR = SpriteTableR_26_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableR = SpriteTableR_26_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableR = SpriteTableR_26_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableR = SpriteTableR_26_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableR = SpriteTableR_26_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableR = SpriteTableR_26_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableR = SpriteTableR_26_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableR = SpriteTableR_26_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableR = SpriteTableR_26_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableR = SpriteTableR_26_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableR = SpriteTableR_26_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableR = SpriteTableR_26_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableR = SpriteTableR_26_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableR = SpriteTableR_26_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableR = SpriteTableR_26_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableR = SpriteTableR_26_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableR = SpriteTableR_26_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableR = SpriteTableR_26_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableR = SpriteTableR_26_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableR = SpriteTableR_27_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableR = SpriteTableR_27_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableR = SpriteTableR_27_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableR = SpriteTableR_27_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableR = SpriteTableR_27_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableR = SpriteTableR_27_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableR = SpriteTableR_27_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableR = SpriteTableR_27_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableR = SpriteTableR_27_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableR = SpriteTableR_27_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableR = SpriteTableR_27_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableR = SpriteTableR_27_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableR = SpriteTableR_27_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_27_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableR = SpriteTableR_27_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableR = SpriteTableR_27_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableR = SpriteTableR_27_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableR = SpriteTableR_27_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableR = SpriteTableR_27_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableR = SpriteTableR_27_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableR = SpriteTableR_27_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableR = SpriteTableR_27_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableR = SpriteTableR_27_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableR = SpriteTableR_27_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableR = SpriteTableR_27_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableR = SpriteTableR_27_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableR = SpriteTableR_27_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableR = SpriteTableR_27_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableR = SpriteTableR_27_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableR = SpriteTableR_27_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableR = SpriteTableR_27_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableR = SpriteTableR_27_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableR = SpriteTableR_27_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableR = SpriteTableR_27_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableR = SpriteTableR_27_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableR = SpriteTableR_27_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableR = SpriteTableR_28_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableR = SpriteTableR_28_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableR = SpriteTableR_28_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableR = SpriteTableR_28_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableR = SpriteTableR_28_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableR = SpriteTableR_28_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableR = SpriteTableR_28_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableR = SpriteTableR_28_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableR = SpriteTableR_28_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableR = SpriteTableR_28_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableR = SpriteTableR_28_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableR = SpriteTableR_28_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableR = SpriteTableR_28_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_28_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableR = SpriteTableR_28_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableR = SpriteTableR_28_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableR = SpriteTableR_28_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableR = SpriteTableR_28_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableR = SpriteTableR_28_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableR = SpriteTableR_28_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableR = SpriteTableR_28_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableR = SpriteTableR_28_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableR = SpriteTableR_28_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableR = SpriteTableR_28_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableR = SpriteTableR_28_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableR = SpriteTableR_28_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableR = SpriteTableR_28_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableR = SpriteTableR_28_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableR = SpriteTableR_28_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableR = SpriteTableR_28_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableR = SpriteTableR_28_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableR = SpriteTableR_28_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableR = SpriteTableR_28_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableR = SpriteTableR_28_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableR = SpriteTableR_28_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableR = SpriteTableR_28_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableR = SpriteTableR_29_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableR = SpriteTableR_29_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableR = SpriteTableR_29_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableR = SpriteTableR_29_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableR = SpriteTableR_29_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableR = SpriteTableR_29_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableR = SpriteTableR_29_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableR = SpriteTableR_29_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableR = SpriteTableR_29_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableR = SpriteTableR_29_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableR = SpriteTableR_29_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableR = SpriteTableR_29_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableR = SpriteTableR_29_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_29_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableR = SpriteTableR_29_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableR = SpriteTableR_29_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableR = SpriteTableR_29_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableR = SpriteTableR_29_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableR = SpriteTableR_29_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableR = SpriteTableR_29_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableR = SpriteTableR_29_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableR = SpriteTableR_29_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableR = SpriteTableR_29_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableR = SpriteTableR_29_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableR = SpriteTableR_29_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableR = SpriteTableR_29_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableR = SpriteTableR_29_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableR = SpriteTableR_29_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableR = SpriteTableR_29_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableR = SpriteTableR_29_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableR = SpriteTableR_29_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableR = SpriteTableR_29_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableR = SpriteTableR_29_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableR = SpriteTableR_29_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableR = SpriteTableR_29_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableR = SpriteTableR_29_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableR = SpriteTableR_30_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableR = SpriteTableR_30_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableR = SpriteTableR_30_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableR = SpriteTableR_30_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableR = SpriteTableR_30_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableR = SpriteTableR_30_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableR = SpriteTableR_30_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableR = SpriteTableR_30_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableR = SpriteTableR_30_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableR = SpriteTableR_30_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableR = SpriteTableR_30_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableR = SpriteTableR_30_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableR = SpriteTableR_30_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_30_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableR = SpriteTableR_30_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableR = SpriteTableR_30_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableR = SpriteTableR_30_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableR = SpriteTableR_30_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableR = SpriteTableR_30_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableR = SpriteTableR_30_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableR = SpriteTableR_30_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableR = SpriteTableR_30_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableR = SpriteTableR_30_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableR = SpriteTableR_30_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableR = SpriteTableR_30_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableR = SpriteTableR_30_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableR = SpriteTableR_30_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableR = SpriteTableR_30_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableR = SpriteTableR_30_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableR = SpriteTableR_30_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableR = SpriteTableR_30_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableR = SpriteTableR_30_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableR = SpriteTableR_30_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableR = SpriteTableR_30_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableR = SpriteTableR_30_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableR = SpriteTableR_30_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableR = SpriteTableR_31_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableR = SpriteTableR_31_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableR = SpriteTableR_31_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableR = SpriteTableR_31_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableR = SpriteTableR_31_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableR = SpriteTableR_31_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableR = SpriteTableR_31_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableR = SpriteTableR_31_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableR = SpriteTableR_31_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableR = SpriteTableR_31_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableR = SpriteTableR_31_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableR = SpriteTableR_31_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableR = SpriteTableR_31_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableR = SpriteTableR_31_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableR = SpriteTableR_31_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableR = SpriteTableR_31_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableR = SpriteTableR_31_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableR = SpriteTableR_31_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableR = SpriteTableR_31_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableR = SpriteTableR_31_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableR = SpriteTableR_31_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableR = SpriteTableR_31_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableR = SpriteTableR_31_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableR = SpriteTableR_31_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableR = SpriteTableR_31_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableR = SpriteTableR_31_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableR = SpriteTableR_31_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableR = SpriteTableR_31_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableR = SpriteTableR_31_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableR = SpriteTableR_31_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableR = SpriteTableR_31_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableR = SpriteTableR_31_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableR = SpriteTableR_31_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableR = SpriteTableR_31_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableR = SpriteTableR_31_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableR = SpriteTableR_31_35[Y_Index][X_Index];
		end
	end

parameter bit [2:0] SpriteTableR_0_0[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_0_1[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_0_2[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_0_3[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_0_4[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_0_5[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_0_6[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd3}};

parameter bit [2:0] SpriteTableR_0_7[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_0_8[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_0_9[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd1,3'd4}};

parameter bit [2:0] SpriteTableR_0_10[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd1,3'd1,3'd1,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd1,3'd1,3'd1,3'd4},
'{3'd4,3'd4,3'd1,3'd1,3'd1,3'd1,3'd1,3'd4},
'{3'd4,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd4},
'{3'd4,3'd1,3'd1,3'd1,3'd1,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_0_11[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_0_12[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_0_13[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_0_14[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_0_15[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_0_16[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_0_17[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_0_18[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_0_19[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_0_20[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_0_21[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_0_22[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_0_23[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_0_24[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_0_25[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_0_26[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2}};

parameter bit [2:0] SpriteTableR_0_27[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_0_28[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_0_29[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_0_30[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_0_31[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_0_32[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_0_33[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_0_34[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1}};

parameter bit [2:0] SpriteTableR_0_35[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_1_0[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_1_1[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_1_2[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_1_3[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_1_4[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_1_5[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd2,3'd3,3'd3,3'd4,3'd1,3'd4},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd3,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_1_6[7:0][7:0] = '{'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_1_7[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_1_8[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd1,3'd4,3'd3,3'd1,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd2,3'd3,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_1_9[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd1,3'd3,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_1_10[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_1_11[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_1_12[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_1_13[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_1_14[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_1_15[7:0][7:0] = '{'{3'd4,3'd1,3'd1,3'd2,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd2,3'd2,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd2,3'd2,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd1,3'd2,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd2,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_1_16[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_1_17[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd2,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd2,3'd1,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd2,3'd2,3'd1,3'd1,3'd4},
'{3'd4,3'd1,3'd1,3'd2,3'd2,3'd1,3'd1,3'd1},
'{3'd4,3'd1,3'd1,3'd2,3'd2,3'd1,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_1_18[7:0][7:0] = '{'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd1,3'd4,3'd2,3'd1,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_1_19[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_1_20[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3}};

parameter bit [2:0] SpriteTableR_1_21[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_1_22[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_1_23[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_1_24[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd2,3'd2,3'd2,3'd1,3'd1,3'd4,3'd4,3'd4},
'{3'd1,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_1_25[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4}};

parameter bit [2:0] SpriteTableR_1_26[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd1,3'd4,3'd4},
'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_1_27[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_1_28[7:0][7:0] = '{'{3'd4,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd2,3'd1,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_1_29[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_1_30[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2}};

parameter bit [2:0] SpriteTableR_1_31[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_1_32[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd1,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_1_33[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_1_34[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1}};

parameter bit [2:0] SpriteTableR_1_35[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_2_0[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_2_1[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_2_2[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_2_3[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_2_4[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_2_5[7:0][7:0] = '{'{3'd4,3'd3,3'd4,3'd4,3'd2,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd2,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4}};

parameter bit [2:0] SpriteTableR_2_6[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3}};

parameter bit [2:0] SpriteTableR_2_7[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd1,3'd4,3'd1,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd3,3'd3,3'd3,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_2_8[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_2_9[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd2,3'd1},
'{3'd4,3'd3,3'd3,3'd3,3'd2,3'd2,3'd1,3'd4},
'{3'd1,3'd1,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_2_10[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_2_11[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_2_12[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd2,3'd4,3'd1,3'd1,3'd1},
'{3'd4,3'd4,3'd1,3'd2,3'd2,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd2,3'd2,3'd2,3'd4,3'd1},
'{3'd4,3'd1,3'd2,3'd2,3'd2,3'd4,3'd4,3'd1},
'{3'd4,3'd1,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_2_13[7:0][7:0] = '{'{3'd4,3'd1,3'd1,3'd1,3'd2,3'd2,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_2_14[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_2_15[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_2_16[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd3,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_2_17[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd1,3'd2,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_2_18[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_2_19[7:0][7:0] = '{'{3'd4,3'd4,3'd1,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_2_20[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_2_21[7:0][7:0] = '{'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd1,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_2_22[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd1,3'd1,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_2_23[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd2,3'd4,3'd2,3'd1,3'd4,3'd4},
'{3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_2_24[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_2_25[7:0][7:0] = '{'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_2_26[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd2,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_2_27[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd1,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_2_28[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd1,3'd4,3'd4,3'd1,3'd1,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd2,3'd2,3'd1},
'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4},
'{3'd4,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4}};

parameter bit [2:0] SpriteTableR_2_29[7:0][7:0] = '{'{3'd4,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd1,3'd2,3'd2,3'd2,3'd2,3'd4},
'{3'd4,3'd4,3'd1,3'd2,3'd2,3'd2,3'd2,3'd4},
'{3'd4,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd1,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4},
'{3'd4,3'd1,3'd1,3'd4,3'd4,3'd1,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd1,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd1,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_2_30[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd2,3'd3,3'd3,3'd1,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_2_31[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_2_32[7:0][7:0] = '{'{3'd2,3'd3,3'd3,3'd1,3'd1,3'd4,3'd3,3'd4},
'{3'd1,3'd4,3'd4,3'd3,3'd3,3'd4,3'd3,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_2_33[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_2_34[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_2_35[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_3_0[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_3_1[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_3_2[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd1,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd1,3'd1,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_3_3[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_3_4[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd1,3'd1},
'{3'd4,3'd4,3'd1,3'd4,3'd3,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_3_5[7:0][7:0] = '{'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_3_6[7:0][7:0] = '{'{3'd3,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd2,3'd1,3'd4,3'd1,3'd3,3'd4,3'd1,3'd4},
'{3'd3,3'd3,3'd4,3'd4,3'd3,3'd1,3'd1,3'd4},
'{3'd3,3'd3,3'd4,3'd4,3'd3,3'd3,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4},
'{3'd3,3'd4,3'd1,3'd4,3'd1,3'd3,3'd4,3'd4},
'{3'd3,3'd3,3'd3,3'd4,3'd4,3'd2,3'd1,3'd4},
'{3'd1,3'd4,3'd3,3'd4,3'd4,3'd2,3'd1,3'd4}};

parameter bit [2:0] SpriteTableR_3_7[7:0][7:0] = '{'{3'd4,3'd3,3'd3,3'd4,3'd4,3'd2,3'd3,3'd4},
'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd1,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd2,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_3_8[7:0][7:0] = '{'{3'd4,3'd4,3'd1,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd1,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd2,3'd2,3'd2,3'd1,3'd1},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd1,3'd1,3'd1},
'{3'd3,3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd4},
'{3'd4,3'd2,3'd1,3'd1,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd1,3'd4,3'd4,3'd1,3'd4,3'd1},
'{3'd1,3'd1,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_3_9[7:0][7:0] = '{'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_3_10[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_3_11[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_3_12[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_3_13[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd3,3'd1,3'd4}};

parameter bit [2:0] SpriteTableR_3_14[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_3_15[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2}};

parameter bit [2:0] SpriteTableR_3_16[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_3_17[7:0][7:0] = '{'{3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2}};

parameter bit [2:0] SpriteTableR_3_18[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd4,3'd4},
'{3'd4,3'd1,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd2,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_3_19[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_3_20[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_3_21[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_3_22[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_3_23[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd1,3'd1},
'{3'd4,3'd4,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_3_24[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd2,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4},
'{3'd3,3'd3,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd4,3'd4,3'd1,3'd4,3'd1,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd2,3'd1,3'd4}};

parameter bit [2:0] SpriteTableR_3_25[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1},
'{3'd1,3'd2,3'd1,3'd1,3'd1,3'd2,3'd2,3'd1},
'{3'd1,3'd2,3'd2,3'd2,3'd2,3'd4,3'd2,3'd1},
'{3'd4,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd4,3'd4,3'd2,3'd2,3'd1,3'd1,3'd1,3'd2},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_3_26[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd1,3'd1,3'd1,3'd4,3'd2,3'd2,3'd4,3'd2},
'{3'd1,3'd1,3'd1,3'd4,3'd4,3'd4,3'd2,3'd2},
'{3'd4,3'd1,3'd4,3'd1,3'd4,3'd2,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd3}};

parameter bit [2:0] SpriteTableR_3_27[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd2,3'd2,3'd1,3'd4,3'd4,3'd3,3'd4,3'd1},
'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_3_28[7:0][7:0] = '{'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_3_29[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd3,3'd4,3'd1,3'd1,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_3_30[7:0][7:0] = '{'{3'd4,3'd1,3'd3,3'd4,3'd3,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd3},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3}};

parameter bit [2:0] SpriteTableR_3_31[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd3}};

parameter bit [2:0] SpriteTableR_3_32[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd3,3'd3,3'd4,3'd4},
'{3'd4,3'd2,3'd3,3'd2,3'd4,3'd1,3'd4,3'd1},
'{3'd1,3'd3,3'd4,3'd3,3'd4,3'd1,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_3_33[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_3_34[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_3_35[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_4_0[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_4_1[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_4_2[7:0][7:0] = '{'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_4_3[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd2,3'd4},
'{3'd4,3'd4,3'd1,3'd1,3'd2,3'd2,3'd2,3'd4}};

parameter bit [2:0] SpriteTableR_4_4[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd4},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd4},
'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd1,3'd3,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd3}};

parameter bit [2:0] SpriteTableR_4_5[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd3,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd3,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_4_6[7:0][7:0] = '{'{3'd4,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd2,3'd3,3'd2},
'{3'd4,3'd4,3'd4,3'd1,3'd2,3'd1,3'd1,3'd1},
'{3'd4,3'd4,3'd1,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_4_7[7:0][7:0] = '{'{3'd2,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_4_8[7:0][7:0] = '{'{3'd2,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd1,3'd4,3'd1,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd4,3'd2,3'd2},
'{3'd4,3'd1,3'd2,3'd1,3'd4,3'd2,3'd2,3'd4},
'{3'd4,3'd1,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd4}};

parameter bit [2:0] SpriteTableR_4_9[7:0][7:0] = '{'{3'd4,3'd4,3'd1,3'd2,3'd2,3'd2,3'd2,3'd4},
'{3'd4,3'd4,3'd1,3'd2,3'd2,3'd2,3'd2,3'd4},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd2,3'd2,3'd1,3'd1,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd1,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_4_10[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd1,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd2,3'd2,3'd2,3'd4},
'{3'd4,3'd4,3'd1,3'd1,3'd2,3'd2,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd2,3'd1}};

parameter bit [2:0] SpriteTableR_4_11[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd1,3'd1,3'd4}};

parameter bit [2:0] SpriteTableR_4_12[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_4_13[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd3,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_4_14[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd3,3'd2,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_4_15[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd1,3'd1,3'd2,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_4_16[7:0][7:0] = '{'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_4_17[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4}};

parameter bit [2:0] SpriteTableR_4_18[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd3,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_4_19[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_4_20[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4}};

parameter bit [2:0] SpriteTableR_4_21[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd3}};

parameter bit [2:0] SpriteTableR_4_22[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_4_23[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd1,3'd1},
'{3'd4,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd1,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd3,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_4_24[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd3,3'd4},
'{3'd1,3'd4,3'd4,3'd1,3'd4,3'd3,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd1,3'd4,3'd3,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd3,3'd4,3'd3},
'{3'd4,3'd1,3'd3,3'd4,3'd4,3'd4,3'd4,3'd3}};

parameter bit [2:0] SpriteTableR_4_25[7:0][7:0] = '{'{3'd1,3'd2,3'd1,3'd4,3'd4,3'd4,3'd1,3'd1},
'{3'd1,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd1,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd1,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd1,3'd2,3'd2,3'd4,3'd4,3'd1,3'd4,3'd1},
'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd2,3'd2,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_4_26[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd2,3'd1,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd4,3'd4,3'd1},
'{3'd2,3'd2,3'd2,3'd4,3'd4,3'd4,3'd3,3'd3},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd3,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd4,3'd3,3'd2,3'd4,3'd1},
'{3'd4,3'd2,3'd1,3'd4,3'd4,3'd1,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_4_27[7:0][7:0] = '{'{3'd4,3'd4,3'd2,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_4_28[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_4_29[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd1,3'd1,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_4_30[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_4_31[7:0][7:0] = '{'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_4_32[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd2,3'd1,3'd4,3'd1,3'd1,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_4_33[7:0][7:0] = '{'{3'd2,3'd1,3'd4,3'd1,3'd1,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_4_34[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_4_35[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_5_0[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_5_1[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_5_2[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_5_3[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_5_4[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd2,3'd1,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd2,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd1,3'd1,3'd4,3'd4,3'd1,3'd4}};

parameter bit [2:0] SpriteTableR_5_5[7:0][7:0] = '{'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd3,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_5_6[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd3,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd3,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_5_7[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_5_8[7:0][7:0] = '{'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd1,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd1,3'd2,3'd2,3'd2,3'd2,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd2,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd2,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd2,3'd4,3'd1,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_5_9[7:0][7:0] = '{'{3'd4,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3}};

parameter bit [2:0] SpriteTableR_5_10[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1},
'{3'd4,3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd1,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_5_11[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_5_12[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_5_13[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_5_14[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_5_15[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_5_16[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_5_17[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd2,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_5_18[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_5_19[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_5_20[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_5_21[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd3,3'd2},
'{3'd4,3'd1,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_5_22[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd2,3'd1,3'd1,3'd1,3'd4}};

parameter bit [2:0] SpriteTableR_5_23[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_5_24[7:0][7:0] = '{'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_5_25[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_5_26[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd3,3'd4,3'd4,3'd1,3'd3},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_5_27[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd1,3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_5_28[7:0][7:0] = '{'{3'd4,3'd1,3'd1,3'd4,3'd4,3'd1,3'd2,3'd2},
'{3'd4,3'd1,3'd2,3'd1,3'd4,3'd2,3'd4,3'd1},
'{3'd1,3'd4,3'd4,3'd2,3'd1,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd1,3'd1,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_5_29[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_5_30[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_5_31[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_5_32[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_5_33[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_5_34[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_5_35[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_6_0[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd1,3'd4,3'd4,3'd1,3'd4}};

parameter bit [2:0] SpriteTableR_6_1[7:0][7:0] = '{'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd1,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_6_2[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_6_3[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd1,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd1,3'd2,3'd2,3'd2,3'd1,3'd1},
'{3'd4,3'd4,3'd1,3'd1,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_6_4[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd2,3'd2,3'd2,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd1,3'd4,3'd4},
'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4}};

parameter bit [2:0] SpriteTableR_6_5[7:0][7:0] = '{'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4},
'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd1,3'd4,3'd1},
'{3'd4,3'd4,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_6_6[7:0][7:0] = '{'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd2}};

parameter bit [2:0] SpriteTableR_6_7[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd1,3'd4,3'd4,3'd1},
'{3'd4,3'd1,3'd4,3'd4,3'd1,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_6_8[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_6_9[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd2,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd1,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd2,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd1,3'd2,3'd4,3'd4,3'd4,3'd3},
'{3'd1,3'd4,3'd2,3'd1,3'd4,3'd4,3'd1,3'd4}};

parameter bit [2:0] SpriteTableR_6_10[7:0][7:0] = '{'{3'd1,3'd4,3'd2,3'd4,3'd4,3'd4,3'd3,3'd4},
'{3'd1,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd3,3'd4,3'd1},
'{3'd2,3'd1,3'd4,3'd4,3'd4,3'd2,3'd2,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd1,3'd1},
'{3'd1,3'd4,3'd4,3'd4,3'd3,3'd2,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd2,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_6_11[7:0][7:0] = '{'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd2,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd2,3'd1,3'd1,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd2,3'd1,3'd1,3'd4,3'd1},
'{3'd4,3'd4,3'd2,3'd2,3'd1,3'd2,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd2,3'd2,3'd2,3'd4,3'd2},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd4,3'd1,3'd1,3'd4,3'd1,3'd1},
'{3'd4,3'd3,3'd4,3'd4,3'd1,3'd2,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_6_12[7:0][7:0] = '{'{3'd4,3'd3,3'd2,3'd1,3'd1,3'd2,3'd4,3'd1},
'{3'd4,3'd4,3'd2,3'd1,3'd4,3'd1,3'd1,3'd1},
'{3'd1,3'd4,3'd2,3'd4,3'd2,3'd2,3'd1,3'd2},
'{3'd4,3'd4,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd3,3'd4,3'd2,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd3,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_6_13[7:0][7:0] = '{'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2},
'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd2,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2},
'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_6_14[7:0][7:0] = '{'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd3,3'd4,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2},
'{3'd3,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd3,3'd4,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd1,3'd4,3'd2,3'd4,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_6_15[7:0][7:0] = '{'{3'd4,3'd4,3'd2,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd3,3'd4,3'd4,3'd2,3'd2,3'd4,3'd2},
'{3'd4,3'd3,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd1,3'd4,3'd2,3'd4,3'd2,3'd4,3'd2},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd1,3'd3,3'd4,3'd2,3'd1,3'd2}};

parameter bit [2:0] SpriteTableR_6_16[7:0][7:0] = '{'{3'd2,3'd4,3'd4,3'd1,3'd4,3'd2,3'd4,3'd1},
'{3'd4,3'd1,3'd4,3'd4,3'd3,3'd4,3'd1,3'd4},
'{3'd4,3'd2,3'd4,3'd4,3'd1,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd3},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_6_17[7:0][7:0] = '{'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_6_18[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_6_19[7:0][7:0] = '{'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_6_20[7:0][7:0] = '{'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd2}};

parameter bit [2:0] SpriteTableR_6_21[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd2,3'd1,3'd2},
'{3'd3,3'd4,3'd4,3'd3,3'd4,3'd2,3'd1,3'd2},
'{3'd4,3'd4,3'd1,3'd3,3'd4,3'd2,3'd2,3'd2},
'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_6_22[7:0][7:0] = '{'{3'd4,3'd4,3'd1,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd3,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd1,3'd2,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd1,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd1,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_6_23[7:0][7:0] = '{'{3'd4,3'd3,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd3,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd3,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd3,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd3,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd3,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd3,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd3,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_6_24[7:0][7:0] = '{'{3'd4,3'd3,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd3,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd3,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd1,3'd3,3'd2,3'd1,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_6_25[7:0][7:0] = '{'{3'd4,3'd4,3'd1,3'd4,3'd2,3'd1,3'd2,3'd2},
'{3'd1,3'd4,3'd4,3'd2,3'd4,3'd2,3'd2,3'd2},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd2},
'{3'd3,3'd1,3'd1,3'd4,3'd2,3'd4,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3}};

parameter bit [2:0] SpriteTableR_6_26[7:0][7:0] = '{'{3'd3,3'd4,3'd4,3'd3,3'd1,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd1,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd3,3'd1,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd3,3'd2,3'd1,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd3},
'{3'd1,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_6_27[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_6_28[7:0][7:0] = '{'{3'd2,3'd2,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_6_29[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_6_30[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd1,3'd1,3'd1,3'd1,3'd4,3'd1},
'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_6_31[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_6_32[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_6_33[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_6_34[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_6_35[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_7_0[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_7_1[7:0][7:0] = '{'{3'd1,3'd1,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_7_2[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_7_3[7:0][7:0] = '{'{3'd2,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_7_4[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_7_5[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd1,3'd3,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd3,3'd4,3'd3,3'd1}};

parameter bit [2:0] SpriteTableR_7_6[7:0][7:0] = '{'{3'd2,3'd1,3'd1,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_7_7[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_7_8[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd1,3'd4,3'd4,3'd1,3'd4,3'd4,3'd1},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd1}};

parameter bit [2:0] SpriteTableR_7_9[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd2,3'd4,3'd1,3'd1,3'd1},
'{3'd4,3'd4,3'd3,3'd4,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd4,3'd2,3'd1,3'd1,3'd2,3'd1},
'{3'd1,3'd4,3'd4,3'd2,3'd1,3'd1,3'd2,3'd1},
'{3'd3,3'd4,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd4,3'd2,3'd1,3'd4,3'd1,3'd1,3'd1,3'd1},
'{3'd4,3'd1,3'd1,3'd2,3'd1,3'd1,3'd2,3'd1},
'{3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1}};

parameter bit [2:0] SpriteTableR_7_10[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd4,3'd2,3'd1,3'd4,3'd2,3'd1},
'{3'd1,3'd1,3'd4,3'd2,3'd1,3'd1,3'd2,3'd1},
'{3'd1,3'd1,3'd4,3'd1,3'd1,3'd1,3'd1,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd4,3'd2,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd4,3'd1,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_7_11[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd4,3'd2,3'd4},
'{3'd1,3'd1,3'd4,3'd1,3'd1,3'd1,3'd2,3'd4},
'{3'd1,3'd1,3'd4,3'd1,3'd1,3'd1,3'd1,3'd4},
'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd1,3'd4,3'd1,3'd1,3'd4,3'd1,3'd2},
'{3'd2,3'd1,3'd1,3'd2,3'd1,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_7_12[7:0][7:0] = '{'{3'd2,3'd1,3'd1,3'd2,3'd1,3'd4,3'd2,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd4,3'd2,3'd4},
'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd2},
'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd3},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd4,3'd4,3'd3},
'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_7_13[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd4,3'd1},
'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd2,3'd4,3'd1},
'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd2,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd2,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd1},
'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd2,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd2,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_7_14[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd2,3'd4,3'd1},
'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd2,3'd4,3'd1},
'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd2,3'd4,3'd1},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd3},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd4,3'd2,3'd4},
'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_7_15[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4},
'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_7_16[7:0][7:0] = '{'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4},
'{3'd1,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd2,3'd2,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd2,3'd1,3'd4,3'd2,3'd2,3'd2},
'{3'd1,3'd3,3'd4,3'd4,3'd4,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd1,3'd3,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_7_17[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_7_18[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4}};

parameter bit [2:0] SpriteTableR_7_19[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd2,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd4,3'd1,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd3,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_7_20[7:0][7:0] = '{'{3'd4,3'd2,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd2},
'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_7_21[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd1},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd1,3'd1},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd4,3'd2,3'd2,3'd2,3'd1,3'd1,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_7_22[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd3},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd3}};

parameter bit [2:0] SpriteTableR_7_23[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd3},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd3},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd3},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd3},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd3},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4}};

parameter bit [2:0] SpriteTableR_7_24[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd1,3'd2,3'd2,3'd2,3'd1,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_7_25[7:0][7:0] = '{'{3'd1,3'd2,3'd2,3'd1,3'd2,3'd2,3'd2,3'd2},
'{3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd1,3'd2,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd1,3'd2,3'd2,3'd1,3'd2,3'd2,3'd2,3'd2},
'{3'd1,3'd2,3'd2,3'd2,3'd1,3'd2,3'd2,3'd2},
'{3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_7_26[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd1,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd1,3'd1,3'd1,3'd1},
'{3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd4,3'd3,3'd2,3'd3,3'd3,3'd3},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd3}};

parameter bit [2:0] SpriteTableR_7_27[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd1,3'd4,3'd4,3'd3,3'd3,3'd1,3'd4},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd3,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_7_28[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd1,3'd4},
'{3'd3,3'd1,3'd4,3'd4,3'd1,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_7_29[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4}};

parameter bit [2:0] SpriteTableR_7_30[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd2,3'd2,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd4,3'd2,3'd2,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_7_31[7:0][7:0] = '{'{3'd4,3'd1,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd1,3'd2,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_7_32[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_7_33[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_7_34[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_7_35[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_8_0[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_8_1[7:0][7:0] = '{'{3'd2,3'd2,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_8_2[7:0][7:0] = '{'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd2,3'd2,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd2,3'd2,3'd2},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd4,3'd1,3'd4,3'd4,3'd2,3'd2,3'd1},
'{3'd2,3'd4,3'd1,3'd1,3'd2,3'd2,3'd1,3'd1}};

parameter bit [2:0] SpriteTableR_8_3[7:0][7:0] = '{'{3'd2,3'd4,3'd4,3'd4,3'd2,3'd1,3'd2,3'd2},
'{3'd2,3'd4,3'd4,3'd4,3'd2,3'd1,3'd1,3'd2},
'{3'd2,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd1,3'd2,3'd1,3'd3,3'd4,3'd1},
'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd3,3'd1,3'd1,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_8_4[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_8_5[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd1},
'{3'd4,3'd1,3'd3,3'd2,3'd4,3'd4,3'd2,3'd3},
'{3'd3,3'd4,3'd2,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_8_6[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_8_7[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2}};

parameter bit [2:0] SpriteTableR_8_8[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd1,3'd1},
'{3'd4,3'd1,3'd4,3'd4,3'd2,3'd1,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd4,3'd4,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd2,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1,3'd2},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd2,3'd1,3'd1,3'd2,3'd1,3'd1,3'd2}};

parameter bit [2:0] SpriteTableR_8_9[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd2,3'd1,3'd1,3'd2,3'd1,3'd1,3'd2},
'{3'd1,3'd2,3'd1,3'd1,3'd2,3'd1,3'd1,3'd2},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd4},
'{3'd1,3'd2,3'd1,3'd1,3'd2,3'd1,3'd4,3'd3},
'{3'd1,3'd4,3'd1,3'd1,3'd1,3'd2,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_8_10[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd4,3'd3,3'd4},
'{3'd1,3'd2,3'd4,3'd1,3'd2,3'd4,3'd4,3'd4},
'{3'd1,3'd2,3'd1,3'd1,3'd4,3'd3,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd1,3'd4,3'd3,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd1,3'd4,3'd3,3'd4,3'd4,3'd1,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4}};

parameter bit [2:0] SpriteTableR_8_11[7:0][7:0] = '{'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd1,3'd4,3'd4,3'd2,3'd3}};

parameter bit [2:0] SpriteTableR_8_12[7:0][7:0] = '{'{3'd3,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd3,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_8_13[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_8_14[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd3,3'd3,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd1,3'd1,3'd4,3'd4,3'd3,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd1,3'd4,3'd4,3'd1,3'd4,3'd4,3'd1},
'{3'd4,3'd2,3'd1,3'd1,3'd3,3'd1,3'd3,3'd4}};

parameter bit [2:0] SpriteTableR_8_15[7:0][7:0] = '{'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd2,3'd4,3'd4,3'd2,3'd2,3'd4},
'{3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd4,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd4,3'd2},
'{3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_8_16[7:0][7:0] = '{'{3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd2,3'd1,3'd4,3'd1,3'd2,3'd2,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd1,3'd4}};

parameter bit [2:0] SpriteTableR_8_17[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd3,3'd4,3'd4,3'd1,3'd1,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd2,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd1,3'd1},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_8_18[7:0][7:0] = '{'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd4,3'd4,3'd2},
'{3'd1,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd1,3'd4,3'd2,3'd1,3'd1,3'd2},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd1,3'd1,3'd1},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2},
'{3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2}};

parameter bit [2:0] SpriteTableR_8_19[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2},
'{3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2},
'{3'd4,3'd2,3'd4,3'd4,3'd2,3'd2,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2}};

parameter bit [2:0] SpriteTableR_8_20[7:0][7:0] = '{'{3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd4,3'd4,3'd3,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd2,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd1},
'{3'd2,3'd2,3'd2,3'd4,3'd1,3'd4,3'd4,3'd3}};

parameter bit [2:0] SpriteTableR_8_21[7:0][7:0] = '{'{3'd2,3'd2,3'd4,3'd3,3'd1,3'd4,3'd1,3'd4},
'{3'd4,3'd2,3'd4,3'd1,3'd4,3'd4,3'd3,3'd4},
'{3'd4,3'd2,3'd2,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd2,3'd4,3'd3,3'd4,3'd4,3'd3,3'd4,3'd4},
'{3'd2,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_8_22[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd3}};

parameter bit [2:0] SpriteTableR_8_23[7:0][7:0] = '{'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd3,3'd1},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd1,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd4,3'd4,3'd1,3'd4,3'd1,3'd3}};

parameter bit [2:0] SpriteTableR_8_24[7:0][7:0] = '{'{3'd4,3'd4,3'd3,3'd3,3'd2,3'd3,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_8_25[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd4,3'd4,3'd2}};

parameter bit [2:0] SpriteTableR_8_26[7:0][7:0] = '{'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd3,3'd1,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd3},
'{3'd4,3'd4,3'd4,3'd1,3'd3,3'd2,3'd4,3'd4},
'{3'd3,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2}};

parameter bit [2:0] SpriteTableR_8_27[7:0][7:0] = '{'{3'd4,3'd1,3'd1,3'd1,3'd1,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd2,3'd4,3'd1},
'{3'd3,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd2,3'd4,3'd1},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd1,3'd4,3'd4,3'd4,3'd3,3'd4}};

parameter bit [2:0] SpriteTableR_8_28[7:0][7:0] = '{'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd2,3'd4,3'd1},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd1,3'd3,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_8_29[7:0][7:0] = '{'{3'd1,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_8_30[7:0][7:0] = '{'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_8_31[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd1,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_8_32[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_8_33[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_8_34[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_8_35[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_9_0[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_9_1[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_9_2[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_9_3[7:0][7:0] = '{'{3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd3,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd2,3'd2,3'd4,3'd3,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd3,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd3,3'd1}};

parameter bit [2:0] SpriteTableR_9_4[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd3,3'd2,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_9_5[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_9_6[7:0][7:0] = '{'{3'd4,3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3}};

parameter bit [2:0] SpriteTableR_9_7[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1},
'{3'd4,3'd4,3'd1,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd2,3'd2,3'd2,3'd1},
'{3'd4,3'd4,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1}};

parameter bit [2:0] SpriteTableR_9_8[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd2,3'd1,3'd1,3'd2,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd2,3'd1,3'd1,3'd2,3'd1,3'd1}};

parameter bit [2:0] SpriteTableR_9_9[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd2,3'd4,3'd4,3'd2,3'd1},
'{3'd1,3'd2,3'd4,3'd4,3'd3,3'd3,3'd4,3'd4},
'{3'd2,3'd4,3'd2,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd1,3'd4,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd1,3'd4}};

parameter bit [2:0] SpriteTableR_9_10[7:0][7:0] = '{'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4},
'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd1,3'd4}};

parameter bit [2:0] SpriteTableR_9_11[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd3,3'd3,3'd4},
'{3'd3,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_9_12[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd2,3'd2},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_9_13[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd2,3'd4,3'd2,3'd4,3'd4,3'd2,3'd2,3'd4},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd3,3'd3,3'd3,3'd1,3'd1,3'd4,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_9_14[7:0][7:0] = '{'{3'd1,3'd4,3'd1,3'd4,3'd3,3'd4,3'd4,3'd2},
'{3'd3,3'd4,3'd1,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd1,3'd4,3'd4,3'd3,3'd4,3'd2,3'd4,3'd1},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd3,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_9_15[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4}};

parameter bit [2:0] SpriteTableR_9_16[7:0][7:0] = '{'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd2,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd1,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_9_17[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4},
'{3'd4,3'd1,3'd3,3'd4,3'd4,3'd4,3'd2,3'd2},
'{3'd4,3'd3,3'd4,3'd2,3'd4,3'd4,3'd1,3'd1},
'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd2,3'd4,3'd2,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd4,3'd1},
'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4}};

parameter bit [2:0] SpriteTableR_9_18[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd4,3'd4,3'd1,3'd1,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd1,3'd1,3'd4},
'{3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd1,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_9_19[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd2,3'd4,3'd4,3'd2,3'd2,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd2,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd3,3'd3},
'{3'd2,3'd4,3'd4,3'd3,3'd1,3'd1,3'd4,3'd4},
'{3'd4,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_9_20[7:0][7:0] = '{'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd1,3'd2,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_9_21[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_9_22[7:0][7:0] = '{'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4}};

parameter bit [2:0] SpriteTableR_9_23[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd2},
'{3'd4,3'd4,3'd1,3'd4,3'd1,3'd2,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd2,3'd2},
'{3'd1,3'd4,3'd4,3'd1,3'd4,3'd2,3'd2,3'd2},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd2,3'd2,3'd2},
'{3'd4,3'd1,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd1,3'd2,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_9_24[7:0][7:0] = '{'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_9_25[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4,3'd3},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd3,3'd4},
'{3'd2,3'd2,3'd2,3'd4,3'd4,3'd3,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_9_26[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd1,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd1,3'd4,3'd1,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_9_27[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd1}};

parameter bit [2:0] SpriteTableR_9_28[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd1,3'd4},
'{3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd3,3'd4,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2}};

parameter bit [2:0] SpriteTableR_9_29[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_9_30[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_9_31[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4}};

parameter bit [2:0] SpriteTableR_9_32[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd4,3'd1,3'd1,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd1,3'd2,3'd1,3'd4}};

parameter bit [2:0] SpriteTableR_9_33[7:0][7:0] = '{'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1},
'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4},
'{3'd4,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4},
'{3'd4,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1},
'{3'd4,3'd2,3'd2,3'd1,3'd1,3'd2,3'd2,3'd1},
'{3'd4,3'd1,3'd1,3'd4,3'd4,3'd1,3'd2,3'd1}};

parameter bit [2:0] SpriteTableR_9_34[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_9_35[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_10_0[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_10_1[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2}};

parameter bit [2:0] SpriteTableR_10_2[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_10_3[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_10_4[7:0][7:0] = '{'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd4,3'd3,3'd1,3'd1,3'd1,3'd1}};

parameter bit [2:0] SpriteTableR_10_5[7:0][7:0] = '{'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd2,3'd3,3'd3,3'd3},
'{3'd4,3'd4,3'd3,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_10_6[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_10_7[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2}};

parameter bit [2:0] SpriteTableR_10_8[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd2,3'd1,3'd1,3'd2,3'd1,3'd1,3'd2,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd2,3'd1,3'd1,3'd2,3'd1,3'd1,3'd2,3'd1}};

parameter bit [2:0] SpriteTableR_10_9[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd4,3'd1,3'd1,3'd2,3'd1,3'd1,3'd2,3'd1},
'{3'd4,3'd2,3'd1,3'd2,3'd1,3'd1,3'd2,3'd1},
'{3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd3,3'd4,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3}};

parameter bit [2:0] SpriteTableR_10_10[7:0][7:0] = '{'{3'd4,3'd3,3'd3,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1},
'{3'd4,3'd4,3'd1,3'd4,3'd3,3'd2,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_10_11[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd3,3'd3,3'd1,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_10_12[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd2,3'd2},
'{3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd2,3'd4},
'{3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4},
'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_10_13[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4},
'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd4,3'd4,3'd2,3'd2,3'd4,3'd2,3'd4},
'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_10_14[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd2,3'd2},
'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd2,3'd2,3'd4,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4,3'd3},
'{3'd2,3'd2,3'd4,3'd2,3'd4,3'd2,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd3,3'd4}};

parameter bit [2:0] SpriteTableR_10_15[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd3,3'd1,3'd4},
'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd1,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd3,3'd4,3'd1,3'd1},
'{3'd2,3'd2,3'd2,3'd4,3'd1,3'd4,3'd4,3'd3},
'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd2,3'd4,3'd3,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd1,3'd3,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4}};

parameter bit [2:0] SpriteTableR_10_16[7:0][7:0] = '{'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd2},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd2,3'd3,3'd4,3'd4,3'd3,3'd4,3'd2},
'{3'd1,3'd4,3'd1,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd3,3'd4,3'd4,3'd1,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_10_17[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd2,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_10_18[7:0][7:0] = '{'{3'd2,3'd4,3'd1,3'd1,3'd4,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd1,3'd1,3'd4,3'd2,3'd1},
'{3'd1,3'd4,3'd4,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4},
'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4}};

parameter bit [2:0] SpriteTableR_10_19[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2},
'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4},
'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd4,3'd2,3'd4},
'{3'd1,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2},
'{3'd4,3'd1,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_10_20[7:0][7:0] = '{'{3'd4,3'd4,3'd2,3'd2,3'd4,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd3,3'd4,3'd1,3'd4,3'd2,3'd2},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd3,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd2,3'd4,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_10_21[7:0][7:0] = '{'{3'd4,3'd4,3'd3,3'd4,3'd2,3'd1,3'd2,3'd2},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd2,3'd4,3'd2,3'd2,3'd2},
'{3'd1,3'd1,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd1,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd3,3'd4,3'd2,3'd4,3'd4,3'd2,3'd2},
'{3'd1,3'd3,3'd4,3'd1,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd2,3'd1,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_10_22[7:0][7:0] = '{'{3'd1,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd3,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_10_23[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd3},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_10_24[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd3,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd2,3'd1,3'd4},
'{3'd2,3'd2,3'd2,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd4,3'd3,3'd4,3'd4,3'd1},
'{3'd2,3'd2,3'd4,3'd2,3'd1,3'd4,3'd4,3'd3},
'{3'd2,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_10_25[7:0][7:0] = '{'{3'd3,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_10_26[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd3,3'd1,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd1,3'd4}};

parameter bit [2:0] SpriteTableR_10_27[7:0][7:0] = '{'{3'd4,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd3,3'd1,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd3,3'd4,3'd3},
'{3'd1,3'd4,3'd4,3'd4,3'd3,3'd4,3'd3,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd1,3'd3,3'd3},
'{3'd4,3'd4,3'd4,3'd1,3'd3,3'd1,3'd3,3'd3}};

parameter bit [2:0] SpriteTableR_10_28[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd3,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd3,3'd1,3'd3,3'd3,3'd1},
'{3'd4,3'd4,3'd1,3'd3,3'd1,3'd3,3'd3,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd3,3'd3,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd3,3'd3,3'd3,3'd4},
'{3'd4,3'd1,3'd3,3'd4,3'd2,3'd3,3'd4,3'd4},
'{3'd4,3'd3,3'd4,3'd1,3'd3,3'd3,3'd1,3'd1},
'{3'd1,3'd3,3'd1,3'd3,3'd3,3'd3,3'd4,3'd3}};

parameter bit [2:0] SpriteTableR_10_29[7:0][7:0] = '{'{3'd4,3'd3,3'd4,3'd3,3'd3,3'd3,3'd4,3'd3},
'{3'd4,3'd3,3'd3,3'd4,3'd4,3'd4,3'd3,3'd4},
'{3'd2,3'd4,3'd2,3'd3,3'd3,3'd2,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_10_30[7:0][7:0] = '{'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_10_31[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_10_32[7:0][7:0] = '{'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd1,3'd4,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd1,3'd1,3'd1,3'd1,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_10_33[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_10_34[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_10_35[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_11_0[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd2,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd1,3'd1,3'd4},
'{3'd1,3'd1,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_11_1[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_11_2[7:0][7:0] = '{'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1},
'{3'd2,3'd2,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1},
'{3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_11_3[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2}};

parameter bit [2:0] SpriteTableR_11_4[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd2},
'{3'd4,3'd1,3'd4,3'd1,3'd4,3'd4,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd1,3'd1,3'd4,3'd1,3'd1,3'd1,3'd1,3'd2}};

parameter bit [2:0] SpriteTableR_11_5[7:0][7:0] = '{'{3'd4,3'd2,3'd1,3'd4,3'd4,3'd1,3'd2,3'd2},
'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd1,3'd4,3'd2},
'{3'd4,3'd1,3'd3,3'd4,3'd2,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd2}};

parameter bit [2:0] SpriteTableR_11_6[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4}};

parameter bit [2:0] SpriteTableR_11_7[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd3,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd3},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_11_8[7:0][7:0] = '{'{3'd1,3'd4,3'd3,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd1,3'd2,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd1,3'd1,3'd2,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd1,3'd1,3'd1,3'd4,3'd3,3'd4,3'd4,3'd4},
'{3'd1,3'd2,3'd1,3'd2,3'd4,3'd4,3'd4,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd4,3'd1,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd4,3'd3,3'd4,3'd4},
'{3'd1,3'd2,3'd1,3'd1,3'd2,3'd2,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_11_9[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd2,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd4,3'd1,3'd4},
'{3'd1,3'd2,3'd1,3'd1,3'd2,3'd4,3'd1,3'd4},
'{3'd1,3'd2,3'd1,3'd1,3'd2,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd3,3'd3,3'd1,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_11_10[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd3,3'd2,3'd3},
'{3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd3,3'd2,3'd3,3'd3,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd1,3'd3,3'd4,3'd1,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_11_11[7:0][7:0] = '{'{3'd3,3'd4,3'd4,3'd4,3'd1,3'd3,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd3,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_11_12[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd2,3'd2,3'd2,3'd4,3'd1,3'd4,3'd3,3'd4},
'{3'd4,3'd2,3'd2,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd4,3'd2,3'd2,3'd4,3'd4,3'd1,3'd4,3'd2},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd3,3'd4,3'd2},
'{3'd4,3'd2,3'd4,3'd3,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd2,3'd4,3'd3,3'd1,3'd4,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_11_13[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd1,3'd3,3'd4,3'd4,3'd2},
'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd2,3'd4,3'd2},
'{3'd4,3'd2,3'd3,3'd4,3'd4,3'd2,3'd4,3'd2},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd2,3'd4,3'd4,3'd3,3'd4,3'd2,3'd2,3'd2},
'{3'd2,3'd4,3'd1,3'd4,3'd2,3'd4,3'd4,3'd2},
'{3'd4,3'd3,3'd1,3'd4,3'd2,3'd4,3'd4,3'd2}};

parameter bit [2:0] SpriteTableR_11_14[7:0][7:0] = '{'{3'd4,3'd3,3'd3,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd3,3'd4,3'd4,3'd2,3'd2,3'd4,3'd4,3'd2},
'{3'd1,3'd4,3'd4,3'd2,3'd2,3'd2,3'd4,3'd2},
'{3'd4,3'd2,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd2,3'd1,3'd2,3'd2,3'd4,3'd2},
'{3'd1,3'd4,3'd2,3'd1,3'd2,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_11_15[7:0][7:0] = '{'{3'd3,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd2,3'd4,3'd4,3'd2,3'd2,3'd4,3'd2},
'{3'd4,3'd2,3'd4,3'd4,3'd2,3'd2,3'd4,3'd2},
'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2},
'{3'd2,3'd2,3'd4,3'd4,3'd2,3'd2,3'd4,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_11_16[7:0][7:0] = '{'{3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd4,3'd4,3'd2},
'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd4,3'd1},
'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_11_17[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd1,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4},
'{3'd4,3'd2,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd2,3'd3,3'd1,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd1,3'd2,3'd3,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_11_18[7:0][7:0] = '{'{3'd1,3'd2,3'd4,3'd1,3'd2,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd1,3'd4,3'd4,3'd3,3'd4},
'{3'd1,3'd2,3'd4,3'd1,3'd1,3'd2,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd2,3'd4,3'd4,3'd2,3'd2,3'd4,3'd3},
'{3'd4,3'd2,3'd4,3'd4,3'd2,3'd2,3'd4,3'd3}};

parameter bit [2:0] SpriteTableR_11_19[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd2,3'd3},
'{3'd4,3'd2,3'd1,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd1,3'd2,3'd4},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd1,3'd2,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd2,3'd3}};

parameter bit [2:0] SpriteTableR_11_20[7:0][7:0] = '{'{3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd2,3'd2},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd2,3'd4},
'{3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd2,3'd3},
'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd2,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd3},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd1},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_11_21[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd4,3'd2,3'd4},
'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4,3'd1},
'{3'd2,3'd2,3'd2,3'd4,3'd2,3'd4,3'd1,3'd1},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd4,3'd4,3'd3,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd3,3'd4,3'd3}};

parameter bit [2:0] SpriteTableR_11_22[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd1,3'd4,3'd1},
'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd4,3'd2,3'd1,3'd4,3'd3},
'{3'd2,3'd2,3'd2,3'd4,3'd3,3'd4,3'd4,3'd1},
'{3'd2,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd3,3'd4,3'd4,3'd4,3'd1},
'{3'd2,3'd2,3'd4,3'd1,3'd4,3'd4,3'd4,3'd3},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3}};

parameter bit [2:0] SpriteTableR_11_23[7:0][7:0] = '{'{3'd2,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd2,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd1,3'd1,3'd4,3'd1,3'd4},
'{3'd1,3'd1,3'd4,3'd3,3'd1,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd1,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_11_24[7:0][7:0] = '{'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd2,3'd4,3'd4,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd3,3'd4},
'{3'd4,3'd4,3'd2,3'd1,3'd4,3'd4,3'd3,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd3,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd1,3'd4,3'd4,3'd2}};

parameter bit [2:0] SpriteTableR_11_25[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd1,3'd4,3'd1},
'{3'd4,3'd3,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd1,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd1,3'd1,3'd4,3'd4,3'd3,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd2}};

parameter bit [2:0] SpriteTableR_11_26[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd2},
'{3'd1,3'd3,3'd1,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd3,3'd1,3'd4,3'd4,3'd3,3'd3,3'd3},
'{3'd4,3'd3,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd3,3'd4,3'd1,3'd3,3'd2,3'd1,3'd4},
'{3'd3,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_11_27[7:0][7:0] = '{'{3'd3,3'd1,3'd4,3'd2,3'd1,3'd1,3'd2,3'd4},
'{3'd3,3'd1,3'd1,3'd1,3'd3,3'd1,3'd1,3'd1},
'{3'd3,3'd1,3'd1,3'd3,3'd4,3'd4,3'd1,3'd1},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd1},
'{3'd1,3'd4,3'd1,3'd1,3'd3,3'd3,3'd1,3'd4},
'{3'd4,3'd3,3'd1,3'd4,3'd1,3'd1,3'd4,3'd4},
'{3'd1,3'd3,3'd4,3'd3,3'd4,3'd4,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_11_28[7:0][7:0] = '{'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd3,3'd1},
'{3'd3,3'd3,3'd4,3'd1,3'd3,3'd3,3'd4,3'd4},
'{3'd3,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd2,3'd3,3'd1,3'd4},
'{3'd4,3'd2,3'd4,3'd3,3'd4,3'd4,3'd3,3'd1},
'{3'd4,3'd2,3'd4,3'd2,3'd4,3'd4,3'd2,3'd1},
'{3'd4,3'd2,3'd4,3'd4,3'd2,3'd2,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_11_29[7:0][7:0] = '{'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd2,3'd2,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4},
'{3'd3,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd1},
'{3'd4,3'd1,3'd4,3'd4,3'd2,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd3,3'd4}};

parameter bit [2:0] SpriteTableR_11_30[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4}};

parameter bit [2:0] SpriteTableR_11_31[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4},
'{3'd1,3'd3,3'd4,3'd3,3'd2,3'd3,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_11_32[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1},
'{3'd4,3'd1,3'd4,3'd4,3'd1,3'd1,3'd1,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd1,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd1,3'd1,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd1,3'd1}};

parameter bit [2:0] SpriteTableR_11_33[7:0][7:0] = '{'{3'd4,3'd4,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1},
'{3'd4,3'd4,3'd1,3'd4,3'd2,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_11_34[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_11_35[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_12_0[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_12_1[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_12_2[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_12_3[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_12_4[7:0][7:0] = '{'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1},
'{3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd2,3'd1},
'{3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd4},
'{3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd4}};

parameter bit [2:0] SpriteTableR_12_5[7:0][7:0] = '{'{3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd4,3'd4},
'{3'd1,3'd2,3'd1,3'd1,3'd1,3'd2,3'd1,3'd4},
'{3'd1,3'd2,3'd1,3'd1,3'd1,3'd2,3'd2,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_12_6[7:0][7:0] = '{'{3'd1,3'd2,3'd4,3'd4,3'd4,3'd2,3'd1,3'd4},
'{3'd1,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd2,3'd1,3'd4,3'd4,3'd2,3'd2,3'd4},
'{3'd2,3'd4,3'd1,3'd4,3'd1,3'd4,3'd4,3'd1},
'{3'd1,3'd3,3'd4,3'd4,3'd4,3'd2,3'd1,3'd4}};

parameter bit [2:0] SpriteTableR_12_7[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd1,3'd4,3'd4,3'd2,3'd2,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd3,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_12_8[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd1,3'd4,3'd2},
'{3'd2,3'd4,3'd2,3'd4,3'd4,3'd1,3'd4,3'd1},
'{3'd3,3'd4,3'd3,3'd4,3'd4,3'd3,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd1}};

parameter bit [2:0] SpriteTableR_12_9[7:0][7:0] = '{'{3'd1,3'd4,3'd1,3'd4,3'd4,3'd4,3'd2,3'd1},
'{3'd1,3'd3,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1},
'{3'd1,3'd4,3'd4,3'd4,3'd3,3'd4,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd1,3'd1},
'{3'd4,3'd4,3'd1,3'd3,3'd4,3'd2,3'd2,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd1,3'd1,3'd1}};

parameter bit [2:0] SpriteTableR_12_10[7:0][7:0] = '{'{3'd4,3'd4,3'd1,3'd4,3'd2,3'd1,3'd1,3'd1},
'{3'd4,3'd4,3'd3,3'd4,3'd1,3'd2,3'd2,3'd1},
'{3'd4,3'd4,3'd3,3'd4,3'd1,3'd2,3'd2,3'd1},
'{3'd4,3'd4,3'd4,3'd2,3'd1,3'd1,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd2,3'd1,3'd2,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd2,3'd4,3'd2,3'd2,3'd4},
'{3'd4,3'd3,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_12_11[7:0][7:0] = '{'{3'd1,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4},
'{3'd3,3'd4,3'd2,3'd4,3'd4,3'd2,3'd2,3'd4},
'{3'd3,3'd2,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4},
'{3'd4,3'd2,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4},
'{3'd4,3'd2,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4}};

parameter bit [2:0] SpriteTableR_12_12[7:0][7:0] = '{'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4}};

parameter bit [2:0] SpriteTableR_12_13[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_12_14[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4}};

parameter bit [2:0] SpriteTableR_12_15[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd2},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd4,3'd4,3'd3},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd2,3'd4,3'd1},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd4,3'd3,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd3,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_12_16[7:0][7:0] = '{'{3'd4,3'd4,3'd2,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd3,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd3,3'd1,3'd4},
'{3'd4,3'd4,3'd2,3'd3,3'd3,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_12_17[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd2,3'd1,3'd1,3'd4,3'd1,3'd1},
'{3'd4,3'd3,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_12_18[7:0][7:0] = '{'{3'd4,3'd3,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd2,3'd1,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd3,3'd2,3'd1,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd3,3'd2,3'd1,3'd1,3'd2,3'd1,3'd4},
'{3'd4,3'd3,3'd2,3'd1,3'd4,3'd4,3'd1,3'd1},
'{3'd4,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd4}};

parameter bit [2:0] SpriteTableR_12_19[7:0][7:0] = '{'{3'd4,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd2,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd1,3'd2,3'd2,3'd1,3'd4,3'd2,3'd2,3'd4},
'{3'd1,3'd2,3'd2,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd1,3'd1,3'd4,3'd4},
'{3'd1,3'd4,3'd2,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd1,3'd4,3'd2,3'd2,3'd4,3'd1,3'd1,3'd4},
'{3'd1,3'd4,3'd2,3'd4,3'd4,3'd4,3'd1,3'd4}};

parameter bit [2:0] SpriteTableR_12_20[7:0][7:0] = '{'{3'd1,3'd4,3'd2,3'd4,3'd4,3'd1,3'd2,3'd4},
'{3'd3,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4},
'{3'd3,3'd4,3'd2,3'd2,3'd4,3'd2,3'd1,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd3,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4}};

parameter bit [2:0] SpriteTableR_12_21[7:0][7:0] = '{'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4},
'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd2,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4},
'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_12_22[7:0][7:0] = '{'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd2,3'd2,3'd2,3'd4,3'd2,3'd2,3'd2},
'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4},
'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1},
'{3'd4,3'd1,3'd2,3'd2,3'd2,3'd1,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_12_23[7:0][7:0] = '{'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd1,3'd4,3'd1},
'{3'd3,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd4,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd1,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd4,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_12_24[7:0][7:0] = '{'{3'd2,3'd2,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd4,3'd1,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd1,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_12_25[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd2}};

parameter bit [2:0] SpriteTableR_12_26[7:0][7:0] = '{'{3'd2,3'd2,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd1,3'd4,3'd1},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd3,3'd3},
'{3'd3,3'd3,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2}};

parameter bit [2:0] SpriteTableR_12_27[7:0][7:0] = '{'{3'd4,3'd2,3'd2,3'd1,3'd1,3'd4,3'd4,3'd4},
'{3'd1,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd1,3'd2,3'd1,3'd4,3'd1,3'd2,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd1,3'd4,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_12_28[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd3},
'{3'd3,3'd2,3'd1,3'd4,3'd1,3'd2,3'd3,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd3},
'{3'd2,3'd2,3'd4,3'd4,3'd1,3'd2,3'd2,3'd1}};

parameter bit [2:0] SpriteTableR_12_29[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd3,3'd1,3'd4,3'd1,3'd3,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd3},
'{3'd3,3'd2,3'd1,3'd4,3'd1,3'd2,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_12_30[7:0][7:0] = '{'{3'd4,3'd4,3'd2,3'd4,3'd3,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd1,3'd4,3'd1,3'd2,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd3,3'd2,3'd1,3'd4,3'd1,3'd2,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_12_31[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd1,3'd4,3'd4,3'd3,3'd3,3'd4},
'{3'd2,3'd4,3'd3,3'd4,3'd1,3'd4,3'd4,3'd1},
'{3'd4,3'd3,3'd1,3'd4,3'd4,3'd3,3'd2,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2},
'{3'd3,3'd4,3'd1,3'd4,3'd1,3'd4,3'd4,3'd2}};

parameter bit [2:0] SpriteTableR_12_32[7:0][7:0] = '{'{3'd1,3'd3,3'd4,3'd4,3'd4,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd1,3'd4,3'd2,3'd2,3'd2,3'd1},
'{3'd1,3'd2,3'd1,3'd2,3'd2,3'd2,3'd1,3'd1},
'{3'd2,3'd2,3'd1,3'd1,3'd2,3'd1,3'd1,3'd2},
'{3'd4,3'd2,3'd2,3'd1,3'd1,3'd2,3'd2,3'd2},
'{3'd1,3'd3,3'd1,3'd2,3'd1,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd1,3'd2,3'd1,3'd1,3'd2},
'{3'd1,3'd1,3'd4,3'd1,3'd2,3'd2,3'd1,3'd1}};

parameter bit [2:0] SpriteTableR_12_33[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd2,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd2,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_12_34[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_12_35[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_13_0[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_13_1[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd1,3'd4,3'd1,3'd1,3'd4,3'd2,3'd2},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd2,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2}};

parameter bit [2:0] SpriteTableR_13_2[7:0][7:0] = '{'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd1},
'{3'd4,3'd1,3'd4,3'd4,3'd2,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd3,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd3,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_13_3[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_13_4[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_13_5[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd3,3'd1,3'd4,3'd4,3'd3,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_13_6[7:0][7:0] = '{'{3'd4,3'd1,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_13_7[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4},
'{3'd3,3'd3,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_13_8[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd2,3'd1,3'd1,3'd2,3'd1,3'd1,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_13_9[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd2,3'd1,3'd1,3'd2,3'd1,3'd1,3'd2,3'd1},
'{3'd2,3'd2,3'd1,3'd2,3'd2,3'd1,3'd2,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2},
'{3'd2,3'd2,3'd1,3'd2,3'd2,3'd1,3'd2,3'd2},
'{3'd1,3'd4,3'd1,3'd1,3'd1,3'd1,3'd1,3'd4}};

parameter bit [2:0] SpriteTableR_13_10[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd4},
'{3'd2,3'd2,3'd1,3'd2,3'd1,3'd1,3'd2,3'd4},
'{3'd2,3'd2,3'd1,3'd2,3'd2,3'd1,3'd2,3'd4},
'{3'd1,3'd1,3'd4,3'd4,3'd1,3'd1,3'd2,3'd4},
'{3'd2,3'd4,3'd4,3'd2,3'd1,3'd1,3'd2,3'd3},
'{3'd2,3'd2,3'd4,3'd2,3'd2,3'd1,3'd4,3'd3},
'{3'd4,3'd4,3'd1,3'd4,3'd1,3'd1,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd2,3'd4}};

parameter bit [2:0] SpriteTableR_13_11[7:0][7:0] = '{'{3'd2,3'd2,3'd4,3'd2,3'd1,3'd1,3'd2,3'd1},
'{3'd2,3'd2,3'd4,3'd2,3'd1,3'd2,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd2,3'd4,3'd1,3'd4},
'{3'd2,3'd2,3'd4,3'd2,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd2,3'd4,3'd1,3'd1,3'd4}};

parameter bit [2:0] SpriteTableR_13_12[7:0][7:0] = '{'{3'd2,3'd2,3'd4,3'd2,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd2,3'd2,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd3,3'd4,3'd1,3'd1},
'{3'd4,3'd4,3'd2,3'd4,3'd1,3'd4,3'd4,3'd1},
'{3'd2,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd2,3'd2,3'd2,3'd4,3'd1,3'd4,3'd1,3'd3},
'{3'd2,3'd2,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_13_13[7:0][7:0] = '{'{3'd4,3'd2,3'd4,3'd1,3'd4,3'd4,3'd4,3'd3},
'{3'd2,3'd2,3'd4,3'd1,3'd4,3'd1,3'd3,3'd2},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd1,3'd2,3'd4,3'd2,3'd4,3'd4,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2},
'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_13_14[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4},
'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4}};

parameter bit [2:0] SpriteTableR_13_15[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd3,3'd3,3'd4,3'd4,3'd2,3'd2},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd1,3'd4,3'd2},
'{3'd4,3'd3,3'd4,3'd1,3'd4,3'd1,3'd4,3'd2},
'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2}};

parameter bit [2:0] SpriteTableR_13_16[7:0][7:0] = '{'{3'd1,3'd4,3'd2,3'd4,3'd4,3'd3,3'd4,3'd4},
'{3'd3,3'd4,3'd3,3'd4,3'd4,3'd3,3'd4,3'd2},
'{3'd3,3'd4,3'd3,3'd4,3'd4,3'd3,3'd4,3'd2},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd3,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd2,3'd4,3'd3},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_13_17[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_13_18[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd2,3'd2,3'd4,3'd2,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd1,3'd4,3'd2,3'd4,3'd2,3'd4,3'd1},
'{3'd1,3'd1,3'd4,3'd2,3'd4,3'd2,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_13_19[7:0][7:0] = '{'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd2,3'd2,3'd2,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd2,3'd4,3'd2,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4},
'{3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd3,3'd4},
'{3'd2,3'd2,3'd4,3'd1,3'd2,3'd4,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_13_20[7:0][7:0] = '{'{3'd1,3'd4,3'd4,3'd2,3'd2,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd4,3'd2,3'd2,3'd4,3'd4,3'd1},
'{3'd2,3'd1,3'd4,3'd4,3'd2,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd2,3'd4,3'd4,3'd1,3'd4},
'{3'd2,3'd2,3'd4,3'd2,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd2,3'd4,3'd3,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_13_21[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd3,3'd1,3'd4},
'{3'd2,3'd2,3'd4,3'd2,3'd4,3'd3,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd2,3'd4,3'd3,3'd4,3'd3},
'{3'd2,3'd2,3'd4,3'd2,3'd4,3'd4,3'd1,3'd4},
'{3'd2,3'd2,3'd4,3'd2,3'd4,3'd1,3'd1,3'd4},
'{3'd2,3'd2,3'd4,3'd2,3'd4,3'd1,3'd4,3'd4},
'{3'd1,3'd1,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd1,3'd2,3'd4,3'd4,3'd3,3'd4}};

parameter bit [2:0] SpriteTableR_13_22[7:0][7:0] = '{'{3'd2,3'd2,3'd4,3'd2,3'd4,3'd4,3'd3,3'd4},
'{3'd2,3'd2,3'd4,3'd2,3'd4,3'd4,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd4,3'd2,3'd4,3'd4,3'd2},
'{3'd2,3'd2,3'd2,3'd4,3'd3,3'd1,3'd4,3'd2},
'{3'd2,3'd2,3'd4,3'd4,3'd3,3'd1,3'd4,3'd2},
'{3'd2,3'd2,3'd2,3'd4,3'd3,3'd3,3'd4,3'd2},
'{3'd2,3'd2,3'd2,3'd4,3'd3,3'd3,3'd4,3'd2},
'{3'd2,3'd2,3'd2,3'd4,3'd4,3'd2,3'd4,3'd2}};

parameter bit [2:0] SpriteTableR_13_23[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd4,3'd4,3'd4,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd4,3'd3,3'd4,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd4,3'd3,3'd4,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd4,3'd3,3'd4,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd4,3'd4,3'd4,3'd2,3'd2},
'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd4,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_13_24[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_13_25[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2}};

parameter bit [2:0] SpriteTableR_13_26[7:0][7:0] = '{'{3'd4,3'd2,3'd3,3'd3,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd1,3'd4,3'd3,3'd3,3'd2,3'd2},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_13_27[7:0][7:0] = '{'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_13_28[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd1,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_13_29[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd2,3'd4,3'd1,3'd1,3'd4}};

parameter bit [2:0] SpriteTableR_13_30[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd2,3'd4},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd1,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd3,3'd4,3'd3,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_13_31[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd2,3'd2},
'{3'd4,3'd2,3'd4,3'd3,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd2,3'd3},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_13_32[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd1,3'd4,3'd4,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd2,3'd4,3'd4,3'd3,3'd3},
'{3'd4,3'd2,3'd2,3'd4,3'd1,3'd4,3'd3,3'd3},
'{3'd2,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_13_33[7:0][7:0] = '{'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd1,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_13_34[7:0][7:0] = '{'{3'd4,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd1},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_13_35[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_14_0[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd2,3'd2},
'{3'd4,3'd4,3'd1,3'd2,3'd4,3'd3,3'd3,3'd3},
'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_14_1[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_14_2[7:0][7:0] = '{'{3'd3,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_14_3[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd1,3'd1,3'd1,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd1,3'd1,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd3,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd3,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd3,3'd2,3'd4}};

parameter bit [2:0] SpriteTableR_14_4[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_14_5[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd3,3'd1,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_14_6[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd1,3'd1,3'd2,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd1,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4}};

parameter bit [2:0] SpriteTableR_14_7[7:0][7:0] = '{'{3'd4,3'd4,3'd1,3'd1,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd1,3'd3},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1},
'{3'd4,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_14_8[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd2,3'd2,3'd1,3'd2,3'd2,3'd1,3'd2}};

parameter bit [2:0] SpriteTableR_14_9[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd2,3'd4,3'd4,3'd1,3'd1,3'd2,3'd1,3'd2},
'{3'd2,3'd4,3'd4,3'd1,3'd2,3'd2,3'd1,3'd2},
'{3'd4,3'd3,3'd4,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd4,3'd3,3'd4,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd4,3'd3,3'd4,3'd1,3'd2,3'd2,3'd1,3'd2},
'{3'd3,3'd3,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1}};

parameter bit [2:0] SpriteTableR_14_10[7:0][7:0] = '{'{3'd3,3'd4,3'd2,3'd1,3'd1,3'd1,3'd4,3'd1},
'{3'd1,3'd3,3'd2,3'd1,3'd1,3'd2,3'd1,3'd2},
'{3'd4,3'd3,3'd2,3'd1,3'd2,3'd2,3'd1,3'd2},
'{3'd4,3'd3,3'd2,3'd1,3'd4,3'd1,3'd1,3'd1},
'{3'd4,3'd3,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1},
'{3'd4,3'd4,3'd1,3'd1,3'd1,3'd2,3'd4,3'd2},
'{3'd4,3'd4,3'd2,3'd1,3'd1,3'd1,3'd1,3'd4},
'{3'd1,3'd4,3'd2,3'd4,3'd1,3'd1,3'd1,3'd4}};

parameter bit [2:0] SpriteTableR_14_11[7:0][7:0] = '{'{3'd1,3'd4,3'd2,3'd4,3'd1,3'd1,3'd1,3'd2},
'{3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd4,3'd2},
'{3'd4,3'd2,3'd1,3'd1,3'd1,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd1,3'd1,3'd2,3'd2,3'd4,3'd2},
'{3'd3,3'd4,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2},
'{3'd3,3'd4,3'd4,3'd4,3'd1,3'd1,3'd1,3'd4},
'{3'd3,3'd2,3'd4,3'd4,3'd1,3'd4,3'd1,3'd4},
'{3'd3,3'd2,3'd2,3'd1,3'd2,3'd2,3'd1,3'd2}};

parameter bit [2:0] SpriteTableR_14_12[7:0][7:0] = '{'{3'd3,3'd2,3'd2,3'd4,3'd2,3'd2,3'd1,3'd2},
'{3'd3,3'd2,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2},
'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2}};

parameter bit [2:0] SpriteTableR_14_13[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2},
'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_14_14[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2},
'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_14_15[7:0][7:0] = '{'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2},
'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_14_16[7:0][7:0] = '{'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd4},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd4},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd4,3'd1},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_14_17[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_14_18[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd2,3'd2,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd1,3'd4,3'd2,3'd4,3'd4,3'd2}};

parameter bit [2:0] SpriteTableR_14_19[7:0][7:0] = '{'{3'd4,3'd4,3'd1,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd3,3'd4,3'd2,3'd2,3'd4,3'd2},
'{3'd4,3'd4,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd2,3'd2,3'd2,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd4,3'd2},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_14_20[7:0][7:0] = '{'{3'd4,3'd3,3'd4,3'd4,3'd2,3'd2,3'd4,3'd2},
'{3'd4,3'd4,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2},
'{3'd4,3'd4,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2},
'{3'd1,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd2,3'd2,3'd4,3'd1},
'{3'd3,3'd4,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2},
'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2}};

parameter bit [2:0] SpriteTableR_14_21[7:0][7:0] = '{'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2},
'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd4,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_14_22[7:0][7:0] = '{'{3'd4,3'd2,3'd1,3'd4,3'd2,3'd2,3'd4,3'd2},
'{3'd4,3'd2,3'd4,3'd1,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_14_23[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd1,3'd2,3'd2,3'd2,3'd1,3'd4},
'{3'd2,3'd2,3'd1,3'd1,3'd2,3'd2,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd4,3'd2,3'd2,3'd2,3'd1},
'{3'd2,3'd2,3'd2,3'd1,3'd2,3'd2,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd2}};

parameter bit [2:0] SpriteTableR_14_24[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd3},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd1},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd1},
'{3'd2,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd4},
'{3'd1,3'd2,3'd2,3'd2,3'd2,3'd4,3'd3,3'd4},
'{3'd1,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4,3'd4},
'{3'd1,3'd2,3'd2,3'd2,3'd2,3'd4,3'd1,3'd4}};

parameter bit [2:0] SpriteTableR_14_25[7:0][7:0] = '{'{3'd2,3'd1,3'd2,3'd1,3'd2,3'd4,3'd1,3'd4},
'{3'd2,3'd2,3'd1,3'd1,3'd2,3'd3,3'd4,3'd4},
'{3'd2,3'd2,3'd1,3'd2,3'd2,3'd3,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd4,3'd4},
'{3'd1,3'd1,3'd2,3'd2,3'd3,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd2,3'd3,3'd1,3'd4,3'd4},
'{3'd3,3'd3,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_14_26[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd1,3'd4,3'd3,3'd3,3'd2,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_14_27[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_14_28[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd3,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd3,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4}};

parameter bit [2:0] SpriteTableR_14_29[7:0][7:0] = '{'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_14_30[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd2,3'd2,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd1,3'd2,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_14_31[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2},
'{3'd4,3'd4,3'd1,3'd1,3'd4,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd3,3'd4,3'd2,3'd2,3'd2,3'd4}};

parameter bit [2:0] SpriteTableR_14_32[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd1,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd1,3'd4,3'd1,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd1,3'd2,3'd1,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_14_33[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_14_34[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_14_35[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_15_0[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd2,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_15_1[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd4,3'd3,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_15_2[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd1,3'd3,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_15_3[7:0][7:0] = '{'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd3,3'd2,3'd3,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd1,3'd3},
'{3'd4,3'd4,3'd4,3'd3,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd2,3'd2,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_15_4[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_15_5[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd1,3'd2,3'd1,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_15_6[7:0][7:0] = '{'{3'd2,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd3,3'd2,3'd4,3'd1},
'{3'd2,3'd1,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd1,3'd4,3'd4,3'd4,3'd1,3'd2},
'{3'd4,3'd2,3'd4,3'd2,3'd2,3'd3,3'd1,3'd2},
'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd2,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd2,3'd2,3'd1,3'd1,3'd2}};

parameter bit [2:0] SpriteTableR_15_7[7:0][7:0] = '{'{3'd4,3'd4,3'd2,3'd4,3'd2,3'd4,3'd2,3'd2},
'{3'd4,3'd4,3'd2,3'd1,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd3},
'{3'd4,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd2,3'd2,3'd1,3'd2,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd4}};

parameter bit [2:0] SpriteTableR_15_8[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd4,3'd2},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd3},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd4,3'd3},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd4,3'd3},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd4,3'd3},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd4,3'd3},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd4,3'd4},
'{3'd2,3'd1,3'd2,3'd2,3'd1,3'd1,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_15_9[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd4,3'd1},
'{3'd2,3'd1,3'd1,3'd2,3'd1,3'd2,3'd4,3'd1},
'{3'd2,3'd1,3'd2,3'd2,3'd1,3'd2,3'd4,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd4,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd4,3'd4},
'{3'd2,3'd1,3'd2,3'd2,3'd1,3'd2,3'd4,3'd4},
'{3'd4,3'd1,3'd1,3'd4,3'd1,3'd2,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_15_10[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd4,3'd4},
'{3'd1,3'd1,3'd2,3'd2,3'd1,3'd2,3'd4,3'd4},
'{3'd1,3'd1,3'd2,3'd2,3'd1,3'd2,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd3,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd3,3'd4},
'{3'd1,3'd1,3'd2,3'd2,3'd1,3'd2,3'd3,3'd4},
'{3'd1,3'd1,3'd4,3'd4,3'd1,3'd2,3'd3,3'd4},
'{3'd1,3'd1,3'd4,3'd4,3'd1,3'd2,3'd3,3'd4}};

parameter bit [2:0] SpriteTableR_15_11[7:0][7:0] = '{'{3'd1,3'd1,3'd2,3'd2,3'd1,3'd2,3'd3,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd4,3'd2,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd4,3'd3,3'd4},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd4,3'd3,3'd4},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd4,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd4,3'd4,3'd4},
'{3'd2,3'd1,3'd1,3'd4,3'd1,3'd4,3'd3,3'd4}};

parameter bit [2:0] SpriteTableR_15_12[7:0][7:0] = '{'{3'd2,3'd1,3'd2,3'd1,3'd1,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd2,3'd4,3'd2,3'd2,3'd2,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd2,3'd2,3'd2,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd2,3'd4,3'd1,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd2,3'd4,3'd1,3'd4},
'{3'd2,3'd4,3'd2,3'd2,3'd2,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd2,3'd2,3'd2,3'd4,3'd1,3'd4}};

parameter bit [2:0] SpriteTableR_15_13[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd2,3'd2,3'd2,3'd4,3'd1,3'd4},
'{3'd2,3'd4,3'd2,3'd2,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd4,3'd4},
'{3'd2,3'd4,3'd2,3'd4,3'd2,3'd2,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd3}};

parameter bit [2:0] SpriteTableR_15_14[7:0][7:0] = '{'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd4,3'd4},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd3,3'd3,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd4},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd3,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd2,3'd4,3'd2},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd4,3'd2,3'd4}};

parameter bit [2:0] SpriteTableR_15_15[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd4,3'd2,3'd2},
'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd4,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd2,3'd2,3'd2},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd4,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_15_16[7:0][7:0] = '{'{3'd2,3'd4,3'd2,3'd4,3'd4,3'd2,3'd2,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd2,3'd4,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd3,3'd3,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_15_17[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd3,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_15_18[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd1,3'd4,3'd2},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_15_19[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd4},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd4,3'd4},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_15_20[7:0][7:0] = '{'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd4,3'd3,3'd4},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd4,3'd3,3'd4},
'{3'd2,3'd4,3'd2,3'd2,3'd2,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd1,3'd4},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd3,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd2,3'd4,3'd1,3'd4,3'd4},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd1,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_15_21[7:0][7:0] = '{'{3'd2,3'd4,3'd2,3'd4,3'd2,3'd4,3'd4,3'd1},
'{3'd2,3'd4,3'd2,3'd4,3'd3,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd2,3'd4,3'd2,3'd4,3'd1,3'd4,3'd1,3'd3},
'{3'd2,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd2,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd3,3'd4,3'd1,3'd3,3'd4}};

parameter bit [2:0] SpriteTableR_15_22[7:0][7:0] = '{'{3'd2,3'd2,3'd4,3'd1,3'd4,3'd4,3'd3,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4},
'{3'd2,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd2},
'{3'd2,3'd4,3'd3,3'd1,3'd4,3'd1,3'd4,3'd2},
'{3'd2,3'd4,3'd1,3'd4,3'd4,3'd1,3'd4,3'd2},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd2},
'{3'd4,3'd2,3'd4,3'd1,3'd4,3'd3,3'd4,3'd2},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd3,3'd4,3'd2}};

parameter bit [2:0] SpriteTableR_15_23[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd1,3'd2},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2},
'{3'd1,3'd4,3'd4,3'd4,3'd1,3'd4,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2},
'{3'd3,3'd4,3'd4,3'd4,3'd3,3'd4,3'd2,3'd2},
'{3'd3,3'd4,3'd1,3'd4,3'd3,3'd4,3'd2,3'd2},
'{3'd1,3'd4,3'd4,3'd4,3'd2,3'd4,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_15_24[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd2,3'd2},
'{3'd1,3'd4,3'd4,3'd4,3'd3,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd2},
'{3'd1,3'd4,3'd1,3'd2,3'd4,3'd2,3'd2,3'd2},
'{3'd1,3'd4,3'd4,3'd2,3'd4,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd3,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd3,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd3,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_15_25[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd1,3'd2},
'{3'd4,3'd4,3'd3,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd3,3'd4,3'd2,3'd1,3'd2,3'd2},
'{3'd4,3'd4,3'd3,3'd4,3'd1,3'd2,3'd2,3'd2},
'{3'd4,3'd1,3'd1,3'd4,3'd1,3'd2,3'd1,3'd2},
'{3'd4,3'd1,3'd3,3'd1,3'd2,3'd2,3'd1,3'd1},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd3,3'd4,3'd2,3'd2,3'd2,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_15_26[7:0][7:0] = '{'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd3,3'd3,3'd4,3'd1,3'd1},
'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd1,3'd1,3'd4,3'd3,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_15_27[7:0][7:0] = '{'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd1,3'd3,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd1,3'd1,3'd4,3'd1,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2},
'{3'd3,3'd3,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_15_28[7:0][7:0] = '{'{3'd4,3'd3,3'd4,3'd1,3'd2,3'd4,3'd2,3'd4},
'{3'd2,3'd4,3'd4,3'd1,3'd4,3'd4,3'd2,3'd2},
'{3'd3,3'd2,3'd3,3'd1,3'd2,3'd2,3'd4,3'd2},
'{3'd3,3'd4,3'd2,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd2,3'd2,3'd4,3'd2,3'd4,3'd1},
'{3'd1,3'd3,3'd2,3'd4,3'd4,3'd4,3'd1,3'd2},
'{3'd1,3'd4,3'd1,3'd4,3'd4,3'd4,3'd1,3'd2},
'{3'd4,3'd4,3'd2,3'd2,3'd4,3'd2,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_15_29[7:0][7:0] = '{'{3'd4,3'd1,3'd2,3'd4,3'd2,3'd2,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd2,3'd4,3'd2,3'd1,3'd4},
'{3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd1,3'd1},
'{3'd1,3'd3,3'd1,3'd4,3'd4,3'd4,3'd1,3'd1},
'{3'd1,3'd1,3'd4,3'd2,3'd4,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd1,3'd3,3'd1,3'd4,3'd4},
'{3'd4,3'd3,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_15_30[7:0][7:0] = '{'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd1,3'd4,3'd3,3'd4,3'd3,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd3,3'd4,3'd3,3'd4,3'd1},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd3,3'd4,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_15_31[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd2,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd2,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd2,3'd1,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd2,3'd4,3'd2,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_15_32[7:0][7:0] = '{'{3'd2,3'd2,3'd4,3'd2,3'd2,3'd2,3'd1,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd1,3'd4,3'd1,3'd2,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_15_33[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_15_34[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_15_35[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_16_0[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_16_1[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd1}};

parameter bit [2:0] SpriteTableR_16_2[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_16_3[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2}};

parameter bit [2:0] SpriteTableR_16_4[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd3,3'd2},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd3,3'd2,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd3,3'd4,3'd3}};

parameter bit [2:0] SpriteTableR_16_5[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd1},
'{3'd3,3'd3,3'd4,3'd4,3'd1,3'd4,3'd2,3'd1},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd3}};

parameter bit [2:0] SpriteTableR_16_6[7:0][7:0] = '{'{3'd2,3'd2,3'd1,3'd4,3'd4,3'd4,3'd3,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd3,3'd4,3'd4,3'd1},
'{3'd3,3'd1,3'd1,3'd4,3'd1,3'd2,3'd3,3'd1},
'{3'd4,3'd1,3'd2,3'd4,3'd1,3'd3,3'd4,3'd1},
'{3'd2,3'd2,3'd2,3'd4,3'd1,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd2,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd1,3'd3,3'd4,3'd2,3'd4}};

parameter bit [2:0] SpriteTableR_16_7[7:0][7:0] = '{'{3'd1,3'd1,3'd4,3'd1,3'd2,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3}};

parameter bit [2:0] SpriteTableR_16_8[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_16_9[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_16_10[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd1,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd2,3'd3,3'd4,3'd4,3'd1,3'd2},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd3,3'd4,3'd1,3'd4,3'd4,3'd3,3'd2},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_16_11[7:0][7:0] = '{'{3'd4,3'd3,3'd3,3'd4,3'd1,3'd1,3'd2,3'd2},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd3,3'd2,3'd1},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd2,3'd2,3'd1},
'{3'd4,3'd3,3'd1,3'd4,3'd1,3'd4,3'd2,3'd2},
'{3'd4,3'd3,3'd4,3'd1,3'd3,3'd4,3'd2,3'd2},
'{3'd4,3'd1,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd1}};

parameter bit [2:0] SpriteTableR_16_12[7:0][7:0] = '{'{3'd4,3'd1,3'd4,3'd3,3'd4,3'd4,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd3,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd2,3'd2},
'{3'd4,3'd4,3'd1,3'd4,3'd2,3'd4,3'd2,3'd2},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd2,3'd4,3'd4,3'd4,3'd2},
'{3'd1,3'd4,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2},
'{3'd4,3'd3,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_16_13[7:0][7:0] = '{'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd2,3'd2,3'd2,3'd4,3'd2,3'd2},
'{3'd3,3'd4,3'd2,3'd2,3'd2,3'd4,3'd2,3'd2},
'{3'd3,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2},
'{3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2},
'{3'd4,3'd2,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2}};

parameter bit [2:0] SpriteTableR_16_14[7:0][7:0] = '{'{3'd2,3'd2,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd1,3'd4,3'd2,3'd4,3'd4,3'd1},
'{3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2},
'{3'd1,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_16_15[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2},
'{3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2},
'{3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_16_16[7:0][7:0] = '{'{3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd4,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd2,3'd2},
'{3'd2,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd2,3'd2,3'd3,3'd3,3'd3},
'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_16_17[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd3,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd2,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd3,3'd3,3'd4,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd1,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd2,3'd3,3'd1,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_16_18[7:0][7:0] = '{'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd2,3'd4,3'd1,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd3,3'd2,3'd4,3'd4,3'd4},
'{3'd2,3'd3,3'd4,3'd4,3'd2,3'd4,3'd2,3'd2},
'{3'd4,3'd3,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd1,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2},
'{3'd2,3'd4,3'd3,3'd4,3'd2,3'd4,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_16_19[7:0][7:0] = '{'{3'd3,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2},
'{3'd4,3'd1,3'd4,3'd2,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2},
'{3'd4,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2},
'{3'd4,3'd3,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_16_20[7:0][7:0] = '{'{3'd4,3'd4,3'd2,3'd4,3'd2,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd4,3'd2,3'd2},
'{3'd4,3'd4,3'd2,3'd4,3'd2,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2},
'{3'd2,3'd4,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2},
'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_16_21[7:0][7:0] = '{'{3'd4,3'd2,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2},
'{3'd4,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2},
'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd4,3'd2,3'd2,3'd2,3'd4,3'd2,3'd2},
'{3'd2,3'd2,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_16_22[7:0][7:0] = '{'{3'd2,3'd2,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd1,3'd4,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_16_23[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd1,3'd1,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd1,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_16_24[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd1,3'd1,3'd2,3'd1,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_16_25[7:0][7:0] = '{'{3'd2,3'd2,3'd1,3'd2,3'd2,3'd2,3'd1,3'd2},
'{3'd2,3'd2,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd1,3'd2,3'd1,3'd1,3'd2},
'{3'd2,3'd2,3'd2,3'd1,3'd2,3'd1,3'd1,3'd2},
'{3'd2,3'd2,3'd1,3'd1,3'd2,3'd2,3'd1,3'd2},
'{3'd2,3'd2,3'd1,3'd2,3'd2,3'd2,3'd1,3'd1},
'{3'd1,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd3}};

parameter bit [2:0] SpriteTableR_16_26[7:0][7:0] = '{'{3'd4,3'd3,3'd3,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1},
'{3'd4,3'd1,3'd4,3'd3,3'd3,3'd2,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd2}};

parameter bit [2:0] SpriteTableR_16_27[7:0][7:0] = '{'{3'd2,3'd4,3'd2,3'd4,3'd2,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd2,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd2,3'd4,3'd2,3'd4,3'd2,3'd1},
'{3'd2,3'd2,3'd4,3'd4,3'd1,3'd2,3'd1,3'd1},
'{3'd4,3'd4,3'd2,3'd2,3'd4,3'd4,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_16_28[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd2,3'd4,3'd2,3'd4,3'd2,3'd4},
'{3'd1,3'd1,3'd1,3'd4,3'd4,3'd2,3'd2,3'd4},
'{3'd4,3'd4,3'd2,3'd1,3'd2,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd2,3'd1,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd2,3'd1,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd1,3'd1,3'd2,3'd4,3'd2,3'd4}};

parameter bit [2:0] SpriteTableR_16_29[7:0][7:0] = '{'{3'd4,3'd4,3'd1,3'd4,3'd1,3'd1,3'd4,3'd4},
'{3'd2,3'd2,3'd1,3'd4,3'd2,3'd4,3'd2,3'd1},
'{3'd4,3'd4,3'd2,3'd1,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd2,3'd1,3'd4,3'd4,3'd4,3'd1},
'{3'd2,3'd2,3'd1,3'd4,3'd2,3'd4,3'd2,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd1},
'{3'd4,3'd3,3'd4,3'd4,3'd1,3'd2,3'd1,3'd1},
'{3'd4,3'd4,3'd3,3'd4,3'd2,3'd4,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_16_30[7:0][7:0] = '{'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd2,3'd4,3'd1,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd3,3'd4,3'd3,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd1,3'd4,3'd4,3'd4,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_16_31[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd2,3'd4,3'd4,3'd1,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd2,3'd4},
'{3'd3,3'd2,3'd4,3'd4,3'd1,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd3,3'd4}};

parameter bit [2:0] SpriteTableR_16_32[7:0][7:0] = '{'{3'd3,3'd3,3'd4,3'd4,3'd1,3'd2,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd1,3'd1,3'd2,3'd4,3'd4},
'{3'd3,3'd2,3'd1,3'd2,3'd2,3'd4,3'd2,3'd4},
'{3'd3,3'd3,3'd4,3'd2,3'd2,3'd2,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd1,3'd4}};

parameter bit [2:0] SpriteTableR_16_33[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_16_34[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_16_35[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_17_0[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_17_1[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_17_2[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_17_3[7:0][7:0] = '{'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd4,3'd2,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd1,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd1,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd2,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd4,3'd2,3'd1,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd2,3'd2,3'd1,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_17_4[7:0][7:0] = '{'{3'd2,3'd2,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd1,3'd4,3'd4,3'd3,3'd1},
'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd2,3'd2,3'd2,3'd1,3'd4,3'd4,3'd1,3'd3},
'{3'd1,3'd4,3'd2,3'd4,3'd4,3'd4,3'd3,3'd4},
'{3'd4,3'd2,3'd2,3'd4,3'd4,3'd4,3'd3,3'd4},
'{3'd4,3'd4,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd3,3'd4,3'd4,3'd3,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_17_5[7:0][7:0] = '{'{3'd3,3'd3,3'd4,3'd4,3'd1,3'd3,3'd4,3'd4},
'{3'd3,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd1,3'd4,3'd4,3'd3,3'd4,3'd1,3'd4},
'{3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd3,3'd2,3'd4,3'd3,3'd4,3'd3,3'd4,3'd3},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd1,3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_17_6[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd3,3'd4,3'd2},
'{3'd1,3'd4,3'd4,3'd3,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd3,3'd2,3'd1,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd3,3'd1},
'{3'd1,3'd4,3'd4,3'd3,3'd4,3'd2,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd2,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_17_7[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd1,3'd3,3'd1,3'd4,3'd1,3'd3,3'd4},
'{3'd1,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd2,3'd4,3'd1,3'd1,3'd4,3'd1,3'd1},
'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd1,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableR_17_8[7:0][7:0] = '{'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd3,3'd4,3'd1,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd2,3'd2,3'd1,3'd1,3'd1},
'{3'd4,3'd4,3'd1,3'd4,3'd2,3'd1,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd1,3'd1,3'd1},
'{3'd4,3'd4,3'd3,3'd4,3'd1,3'd1,3'd1,3'd1},
'{3'd4,3'd4,3'd3,3'd2,3'd1,3'd1,3'd1,3'd1},
'{3'd4,3'd1,3'd4,3'd2,3'd1,3'd2,3'd1,3'd1}};

parameter bit [2:0] SpriteTableR_17_9[7:0][7:0] = '{'{3'd4,3'd1,3'd4,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd4,3'd3,3'd4,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd4,3'd3,3'd4,3'd1,3'd1,3'd2,3'd1,3'd1},
'{3'd4,3'd4,3'd2,3'd1,3'd1,3'd2,3'd1,3'd1},
'{3'd1,3'd4,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd3,3'd4,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd3,3'd4,3'd2,3'd1,3'd2,3'd2,3'd1,3'd2},
'{3'd4,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd4}};

parameter bit [2:0] SpriteTableR_17_10[7:0][7:0] = '{'{3'd4,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd4,3'd2,3'd2,3'd4,3'd1,3'd1,3'd1,3'd2},
'{3'd2,3'd1,3'd2,3'd4,3'd1,3'd1,3'd1,3'd4},
'{3'd1,3'd1,3'd1,3'd4,3'd1,3'd1,3'd1,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd1,3'd1,3'd1},
'{3'd1,3'd4,3'd4,3'd4,3'd1,3'd1,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_17_11[7:0][7:0] = '{'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1,3'd2},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd4},
'{3'd1,3'd2,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd4,3'd1,3'd1,3'd4,3'd1,3'd4},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd1,3'd1}};

parameter bit [2:0] SpriteTableR_17_12[7:0][7:0] = '{'{3'd4,3'd1,3'd2,3'd4,3'd1,3'd2,3'd1,3'd2},
'{3'd1,3'd4,3'd1,3'd1,3'd1,3'd4,3'd4,3'd2},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd2,3'd4},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd2,3'd4}};

parameter bit [2:0] SpriteTableR_17_13[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd3},
'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd3,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd3,3'd1},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd2,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_17_14[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd4,3'd4,3'd3,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd2,3'd4,3'd1,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd2,3'd2,3'd3,3'd1,3'd4,3'd1},
'{3'd4,3'd2,3'd2,3'd4,3'd3,3'd1,3'd4,3'd3},
'{3'd4,3'd4,3'd2,3'd4,3'd1,3'd4,3'd4,3'd3},
'{3'd2,3'd2,3'd2,3'd4,3'd4,3'd1,3'd4,3'd3}};

parameter bit [2:0] SpriteTableR_17_15[7:0][7:0] = '{'{3'd2,3'd2,3'd4,3'd3,3'd4,3'd1,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd2,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd3,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4}};

parameter bit [2:0] SpriteTableR_17_16[7:0][7:0] = '{'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd1,3'd3},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_17_17[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd4,3'd4,3'd3,3'd3,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_17_18[7:0][7:0] = '{'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_17_19[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd4},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4}};

parameter bit [2:0] SpriteTableR_17_20[7:0][7:0] = '{'{3'd4,3'd2,3'd2,3'd4,3'd4,3'd2,3'd2,3'd4},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd3},
'{3'd4,3'd2,3'd2,3'd4,3'd4,3'd2,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd1},
'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_17_21[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd2},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_17_22[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd2,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd2,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd3,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd1,3'd4,3'd1},
'{3'd2,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd4,3'd3,3'd4,3'd4,3'd3}};

parameter bit [2:0] SpriteTableR_17_23[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd4,3'd3,3'd4,3'd4,3'd3},
'{3'd2,3'd2,3'd2,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd2,3'd2,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd3,3'd4,3'd4,3'd3,3'd4},
'{3'd2,3'd2,3'd4,3'd3,3'd4,3'd4,3'd4,3'd3},
'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_17_24[7:0][7:0] = '{'{3'd2,3'd2,3'd4,3'd1,3'd1,3'd4,3'd4,3'd1},
'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4},
'{3'd2,3'd2,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd1,3'd2,3'd2,3'd1,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd2,3'd2},
'{3'd1,3'd1,3'd2,3'd2,3'd2,3'd1,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_17_25[7:0][7:0] = '{'{3'd2,3'd2,3'd1,3'd2,3'd2,3'd1,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd1},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd2,3'd1},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd2,3'd2},
'{3'd1,3'd1,3'd1,3'd2,3'd4,3'd2,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd2,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_17_26[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd3},
'{3'd4,3'd3,3'd3,3'd3,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_17_27[7:0][7:0] = '{'{3'd4,3'd2,3'd4,3'd2,3'd2,3'd2,3'd4,3'd3},
'{3'd4,3'd2,3'd2,3'd2,3'd1,3'd2,3'd4,3'd3},
'{3'd2,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd1,3'd2,3'd4,3'd1,3'd1,3'd2,3'd4,3'd2},
'{3'd4,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_17_28[7:0][7:0] = '{'{3'd2,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd1,3'd4,3'd2,3'd4,3'd2},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd2,3'd4,3'd4,3'd1,3'd4,3'd2,3'd4,3'd2},
'{3'd2,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd2,3'd1,3'd2,3'd4,3'd2}};

parameter bit [2:0] SpriteTableR_17_29[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd2,3'd2,3'd1,3'd4,3'd1,3'd2,3'd1},
'{3'd1,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd2,3'd2,3'd1,3'd4,3'd1,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd1,3'd4,3'd4,3'd3,3'd4,3'd3,3'd4,3'd2}};

parameter bit [2:0] SpriteTableR_17_30[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd3,3'd2,3'd1,3'd4,3'd4,3'd2,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd1,3'd4,3'd1,3'd4,3'd1},
'{3'd1,3'd4,3'd4,3'd3,3'd4,3'd3,3'd4,3'd2},
'{3'd4,3'd3,3'd2,3'd1,3'd4,3'd1,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_17_31[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd3,3'd4,3'd4,3'd1,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd3,3'd3,3'd4,3'd4,3'd1,3'd3,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_17_32[7:0][7:0] = '{'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd3,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd3,3'd4,3'd4,3'd4,3'd3,3'd1},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_17_33[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_17_34[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_17_35[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_18_0[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_18_1[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_18_2[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd2,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd2,3'd2,3'd4,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_18_3[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd4,3'd1},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd1,3'd2,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd1,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_18_4[7:0][7:0] = '{'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd3,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd3},
'{3'd1,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd1,3'd4}};

parameter bit [2:0] SpriteTableR_18_5[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd1,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3}};

parameter bit [2:0] SpriteTableR_18_6[7:0][7:0] = '{'{3'd4,3'd1,3'd4,3'd4,3'd3,3'd4,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4},
'{3'd1,3'd3,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd3,3'd4,3'd3,3'd2}};

parameter bit [2:0] SpriteTableR_18_7[7:0][7:0] = '{'{3'd4,3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd3,3'd3,3'd1,3'd4,3'd4,3'd4},
'{3'd1,3'd3,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd3,3'd3,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4},
'{3'd3,3'd3,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_18_8[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd2,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd2,3'd1,3'd1,3'd2,3'd1,3'd1,3'd2,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd2,3'd1,3'd1,3'd2,3'd1,3'd1,3'd2,3'd1}};

parameter bit [2:0] SpriteTableR_18_9[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd2,3'd1,3'd1,3'd2,3'd1,3'd1,3'd2,3'd1},
'{3'd2,3'd1,3'd1,3'd2,3'd1,3'd1,3'd2,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd2,3'd1,3'd2,3'd2,3'd1,3'd4,3'd2,3'd1},
'{3'd4,3'd1,3'd1,3'd4,3'd1,3'd1,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_18_10[7:0][7:0] = '{'{3'd1,3'd4,3'd1,3'd1,3'd4,3'd1,3'd1,3'd1},
'{3'd2,3'd1,3'd4,3'd2,3'd1,3'd4,3'd2,3'd4},
'{3'd2,3'd1,3'd4,3'd2,3'd1,3'd4,3'd2,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd4,3'd4,3'd1,3'd4},
'{3'd1,3'd1,3'd1,3'd2,3'd4,3'd4,3'd2,3'd4},
'{3'd1,3'd1,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_18_11[7:0][7:0] = '{'{3'd1,3'd1,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4},
'{3'd1,3'd1,3'd1,3'd2,3'd4,3'd4,3'd2,3'd4},
'{3'd4,3'd1,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4}};

parameter bit [2:0] SpriteTableR_18_12[7:0][7:0] = '{'{3'd4,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4},
'{3'd4,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4},
'{3'd3,3'd4,3'd2,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd3,3'd4,3'd2,3'd2,3'd4,3'd4,3'd2,3'd4},
'{3'd3,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd2},
'{3'd3,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4}};

parameter bit [2:0] SpriteTableR_18_13[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd3,3'd2,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4},
'{3'd2,3'd2,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4},
'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd2,3'd4,3'd2,3'd4,3'd2,3'd2,3'd4},
'{3'd4,3'd2,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4}};

parameter bit [2:0] SpriteTableR_18_14[7:0][7:0] = '{'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4},
'{3'd1,3'd4,3'd4,3'd1,3'd1,3'd1,3'd2,3'd4},
'{3'd1,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_18_15[7:0][7:0] = '{'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4},
'{3'd2,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd4,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_18_16[7:0][7:0] = '{'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd1},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd1},
'{3'd2,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd1,3'd1,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_18_17[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd1,3'd1,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_18_18[7:0][7:0] = '{'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd1},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd1,3'd1,3'd1,3'd1,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_18_19[7:0][7:0] = '{'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_18_20[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd1,3'd4,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_18_21[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd4,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd2,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_18_22[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3}};

parameter bit [2:0] SpriteTableR_18_23[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_18_24[7:0][7:0] = '{'{3'd3,3'd4,3'd1,3'd3,3'd4,3'd3,3'd2,3'd4},
'{3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd3,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd3,3'd1},
'{3'd2,3'd1,3'd2,3'd2,3'd2,3'd4,3'd2,3'd4}};

parameter bit [2:0] SpriteTableR_18_25[7:0][7:0] = '{'{3'd1,3'd1,3'd2,3'd2,3'd2,3'd4,3'd3,3'd3},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4,3'd3},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd3,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd3,3'd3,3'd3,3'd4,3'd1,3'd3,3'd2},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4}};

parameter bit [2:0] SpriteTableR_18_26[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd3,3'd4,3'd4,3'd1,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd3,3'd3,3'd2,3'd4,3'd4,3'd2},
'{3'd3,3'd3,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4}};

parameter bit [2:0] SpriteTableR_18_27[7:0][7:0] = '{'{3'd4,3'd4,3'd2,3'd2,3'd1,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd2,3'd2,3'd1,3'd4,3'd1,3'd4},
'{3'd1,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd1,3'd2,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd2,3'd1,3'd4,3'd1,3'd2},
'{3'd4,3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd1},
'{3'd1,3'd1,3'd4,3'd4,3'd2,3'd4,3'd2,3'd4}};

parameter bit [2:0] SpriteTableR_18_28[7:0][7:0] = '{'{3'd1,3'd2,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd2,3'd4,3'd1,3'd4,3'd1,3'd2},
'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd4,3'd4,3'd1,3'd4,3'd1,3'd4},
'{3'd1,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd1,3'd4,3'd1,3'd2}};

parameter bit [2:0] SpriteTableR_18_29[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd2,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd1,3'd4,3'd4,3'd2,3'd4,3'd3,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd3,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd2,3'd2,3'd4,3'd4,3'd1,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_18_30[7:0][7:0] = '{'{3'd1,3'd1,3'd4,3'd4,3'd3,3'd4,3'd3,3'd4},
'{3'd4,3'd4,3'd1,3'd3,3'd1,3'd4,3'd1,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd3,3'd2,3'd1,3'd4,3'd1,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_18_31[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd1,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd3,3'd2,3'd4,3'd4,3'd4,3'd3}};

parameter bit [2:0] SpriteTableR_18_32[7:0][7:0] = '{'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_18_33[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd1,3'd1,3'd4,3'd4,3'd1,3'd4},
'{3'd2,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_18_34[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd1,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_18_35[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_19_0[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_19_1[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_19_2[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd1,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd4,3'd4,3'd4},
'{3'd1,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd2,3'd2,3'd1,3'd1,3'd4,3'd4},
'{3'd1,3'd2,3'd2,3'd1,3'd1,3'd1,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_19_3[7:0][7:0] = '{'{3'd4,3'd2,3'd1,3'd1,3'd2,3'd1,3'd4,3'd4},
'{3'd2,3'd2,3'd1,3'd1,3'd2,3'd2,3'd1,3'd4},
'{3'd1,3'd2,3'd2,3'd1,3'd1,3'd2,3'd2,3'd1},
'{3'd1,3'd2,3'd2,3'd2,3'd1,3'd1,3'd2,3'd2},
'{3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd2},
'{3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd4},
'{3'd1,3'd2,3'd2,3'd2,3'd4,3'd1,3'd4,3'd4},
'{3'd1,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_19_4[7:0][7:0] = '{'{3'd1,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd1,3'd1,3'd3,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd4},
'{3'd4,3'd1,3'd1,3'd1,3'd1,3'd1,3'd4,3'd4},
'{3'd3,3'd4,3'd1,3'd2,3'd4,3'd1,3'd4,3'd1},
'{3'd3,3'd4,3'd1,3'd2,3'd4,3'd1,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_19_5[7:0][7:0] = '{'{3'd4,3'd4,3'd1,3'd1,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd1,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd1,3'd2,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd1,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd1,3'd2,3'd1,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd1,3'd1,3'd1,3'd1,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_19_6[7:0][7:0] = '{'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd1,3'd1,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd2,3'd1,3'd1,3'd2,3'd1,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_19_7[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd3,3'd3,3'd3,3'd2,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_19_8[7:0][7:0] = '{'{3'd1,3'd2,3'd1,3'd1,3'd1,3'd2,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd3,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd4,3'd3,3'd4},
'{3'd1,3'd2,3'd1,3'd1,3'd2,3'd4,3'd3,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd2,3'd4,3'd1,3'd4},
'{3'd1,3'd2,3'd1,3'd1,3'd2,3'd4,3'd1,3'd4}};

parameter bit [2:0] SpriteTableR_19_9[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd2,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd4,3'd4},
'{3'd1,3'd2,3'd1,3'd1,3'd4,3'd3,3'd4,3'd4},
'{3'd1,3'd2,3'd1,3'd1,3'd4,3'd3,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd4,3'd3,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd1,3'd2,3'd4,3'd1,3'd4,3'd1},
'{3'd1,3'd4,3'd1,3'd2,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_19_10[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd1,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd1,3'd2,3'd3,3'd4,3'd4,3'd3},
'{3'd1,3'd4,3'd1,3'd4,3'd3,3'd4,3'd4,3'd3},
'{3'd4,3'd2,3'd4,3'd4,3'd3,3'd4,3'd1,3'd4},
'{3'd4,3'd2,3'd2,3'd4,3'd3,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd1,3'd4,3'd3,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd2}};

parameter bit [2:0] SpriteTableR_19_11[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd2,3'd2,3'd2,3'd1,3'd3,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd2,3'd4},
'{3'd4,3'd2,3'd4,3'd3,3'd4,3'd4,3'd2,3'd2},
'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2},
'{3'd4,3'd2,3'd4,3'd1,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd3,3'd4,3'd4,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_19_12[7:0][7:0] = '{'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd3,3'd3,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd4,3'd4,3'd2},
'{3'd2,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd2,3'd4,3'd4,3'd2,3'd1,3'd1,3'd2}};

parameter bit [2:0] SpriteTableR_19_13[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd2,3'd2,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_19_14[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4},
'{3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd2,3'd2,3'd4,3'd1},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd2,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd1,3'd4},
'{3'd2,3'd2,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_19_15[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd2,3'd4,3'd1,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd4,3'd2,3'd1,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd3,3'd1,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_19_16[7:0][7:0] = '{'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd3,3'd1,3'd4},
'{3'd3,3'd4,3'd1,3'd4,3'd4,3'd2,3'd1,3'd4},
'{3'd2,3'd3,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_19_17[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd1,3'd4},
'{3'd3,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd2,3'd2,3'd1,3'd1,3'd1,3'd2},
'{3'd1,3'd4,3'd4,3'd1,3'd1,3'd4,3'd1,3'd2},
'{3'd4,3'd4,3'd1,3'd1,3'd4,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd1,3'd1,3'd4,3'd4,3'd2,3'd2},
'{3'd1,3'd4,3'd4,3'd1,3'd1,3'd4,3'd4,3'd3},
'{3'd1,3'd4,3'd4,3'd4,3'd1,3'd1,3'd2,3'd4}};

parameter bit [2:0] SpriteTableR_19_18[7:0][7:0] = '{'{3'd1,3'd2,3'd4,3'd4,3'd2,3'd4,3'd2,3'd1},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd4},
'{3'd1,3'd2,3'd1,3'd1,3'd1,3'd2,3'd3,3'd1},
'{3'd1,3'd2,3'd2,3'd1,3'd1,3'd2,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd1,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3}};

parameter bit [2:0] SpriteTableR_19_19[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd1,3'd2},
'{3'd2,3'd1,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_19_20[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd1,3'd4,3'd4,3'd1,3'd3,3'd4,3'd2},
'{3'd4,3'd3,3'd1,3'd4,3'd1,3'd3,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd4},
'{3'd2,3'd4,3'd1,3'd4,3'd1,3'd4,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_19_21[7:0][7:0] = '{'{3'd2,3'd4,3'd1,3'd4,3'd3,3'd4,3'd2,3'd2},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2},
'{3'd2,3'd4,3'd4,3'd4,3'd3,3'd4,3'd2,3'd2},
'{3'd2,3'd4,3'd4,3'd4,3'd2,3'd4,3'd2,3'd2},
'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd2,3'd2,3'd2},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd2,3'd4,3'd2},
'{3'd4,3'd3,3'd4,3'd1,3'd4,3'd2,3'd2,3'd2},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_19_22[7:0][7:0] = '{'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd2,3'd2,3'd2},
'{3'd2,3'd4,3'd4,3'd3,3'd4,3'd4,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd2,3'd2},
'{3'd4,3'd4,3'd1,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd1,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd3,3'd4,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_19_23[7:0][7:0] = '{'{3'd4,3'd4,3'd3,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd1,3'd4,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd1,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd1,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd1,3'd3,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd1,3'd2,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd2,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd1,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_19_24[7:0][7:0] = '{'{3'd1,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd3,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd3,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_19_25[7:0][7:0] = '{'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3}};

parameter bit [2:0] SpriteTableR_19_26[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd3,3'd4,3'd4},
'{3'd1,3'd3,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4}};

parameter bit [2:0] SpriteTableR_19_27[7:0][7:0] = '{'{3'd2,3'd1,3'd4,3'd1,3'd4,3'd4,3'd1,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd3,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd3,3'd2,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd1,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd1,3'd4,3'd4,3'd3,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_19_28[7:0][7:0] = '{'{3'd4,3'd3,3'd3,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd1,3'd4,3'd4,3'd1,3'd2,3'd1,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd1,3'd1,3'd4,3'd4,3'd2,3'd4,3'd2},
'{3'd2,3'd4,3'd4,3'd1,3'd2,3'd1,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_19_29[7:0][7:0] = '{'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd1,3'd4,3'd3,3'd1,3'd4,3'd4},
'{3'd4,3'd1,3'd1,3'd4,3'd4,3'd3,3'd4,3'd3},
'{3'd4,3'd1,3'd1,3'd4,3'd4,3'd3,3'd4,3'd3},
'{3'd3,3'd4,3'd4,3'd4,3'd3,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd2,3'd1,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_19_30[7:0][7:0] = '{'{3'd4,3'd2,3'd2,3'd4,3'd4,3'd1,3'd4,3'd1},
'{3'd1,3'd4,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1},
'{3'd4,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4},
'{3'd4,3'd4,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd4},
'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd2,3'd2,3'd2},
'{3'd1,3'd4,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_19_31[7:0][7:0] = '{'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd2,3'd2,3'd2},
'{3'd1,3'd1,3'd1,3'd4,3'd4,3'd4,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_19_32[7:0][7:0] = '{'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_19_33[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_19_34[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_19_35[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_20_0[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_20_1[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_20_2[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_20_3[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_20_4[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd4},
'{3'd3,3'd1,3'd4,3'd4,3'd1,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd2,3'd1,3'd1,3'd2,3'd4,3'd1,3'd4},
'{3'd4,3'd2,3'd1,3'd1,3'd2,3'd4,3'd1,3'd4}};

parameter bit [2:0] SpriteTableR_20_5[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd1,3'd1,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_20_6[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_20_7[7:0][7:0] = '{'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd1,3'd4,3'd4,3'd1},
'{3'd4,3'd1,3'd4,3'd3,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4}};

parameter bit [2:0] SpriteTableR_20_8[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd2},
'{3'd4,3'd3,3'd3,3'd4,3'd4,3'd3,3'd4,3'd1},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd2,3'd2,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd2,3'd1},
'{3'd4,3'd1,3'd4,3'd4,3'd3,3'd4,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd2,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd2,3'd1,3'd1}};

parameter bit [2:0] SpriteTableR_20_9[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd1,3'd1,3'd1},
'{3'd4,3'd4,3'd1,3'd4,3'd1,3'd1,3'd1,3'd1},
'{3'd4,3'd4,3'd3,3'd4,3'd1,3'd2,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd2,3'd1,3'd2,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd4,3'd3,3'd4,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd4,3'd4,3'd2,3'd1,3'd1,3'd2,3'd1,3'd1},
'{3'd4,3'd4,3'd2,3'd1,3'd1,3'd4,3'd1,3'd1}};

parameter bit [2:0] SpriteTableR_20_10[7:0][7:0] = '{'{3'd3,3'd4,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd4,3'd2,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd2,3'd2,3'd4,3'd1,3'd2,3'd4,3'd1},
'{3'd4,3'd1,3'd1,3'd4,3'd4,3'd1,3'd4,3'd1},
'{3'd2,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_20_11[7:0][7:0] = '{'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd2}};

parameter bit [2:0] SpriteTableR_20_12[7:0][7:0] = '{'{3'd4,3'd4,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd2,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd2,3'd2,3'd4,3'd4},
'{3'd2,3'd4,3'd2,3'd3,3'd4,3'd4,3'd1,3'd2},
'{3'd4,3'd4,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd3,3'd4,3'd1,3'd4,3'd2},
'{3'd4,3'd2,3'd4,3'd3,3'd4,3'd2,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_20_13[7:0][7:0] = '{'{3'd4,3'd4,3'd3,3'd3,3'd2,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd3,3'd4,3'd2,3'd2,3'd2,3'd4},
'{3'd2,3'd4,3'd3,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd3,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd2,3'd2,3'd4,3'd4},
'{3'd4,3'd1,3'd3,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd3,3'd4,3'd3,3'd4,3'd2,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd2,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_20_14[7:0][7:0] = '{'{3'd1,3'd4,3'd2,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd1,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd3,3'd2,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd2,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd1,3'd4,3'd2,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd2,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_20_15[7:0][7:0] = '{'{3'd4,3'd3,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd3,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd3,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd3,3'd4,3'd4,3'd2,3'd2,3'd4,3'd2},
'{3'd4,3'd2,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_20_16[7:0][7:0] = '{'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd1,3'd1,3'd1},
'{3'd1,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd1,3'd4,3'd2,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd3,3'd3,3'd4,3'd1,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd1,3'd1}};

parameter bit [2:0] SpriteTableR_20_17[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd1,3'd4,3'd4,3'd1,3'd4,3'd2,3'd4,3'd4},
'{3'd1,3'd3,3'd2,3'd3,3'd4,3'd4,3'd2,3'd2},
'{3'd4,3'd4,3'd2,3'd1,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd1,3'd1,3'd1,3'd1,3'd4,3'd4},
'{3'd3,3'd2,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_20_18[7:0][7:0] = '{'{3'd3,3'd2,3'd4,3'd1,3'd4,3'd2,3'd4,3'd1},
'{3'd3,3'd2,3'd4,3'd1,3'd4,3'd4,3'd4,3'd1},
'{3'd2,3'd2,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd2,3'd1,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd1,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd2,3'd4,3'd2,3'd4,3'd4,3'd1,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_20_19[7:0][7:0] = '{'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd2,3'd4,3'd4,3'd1,3'd4,3'd1},
'{3'd2,3'd4,3'd2,3'd4,3'd1,3'd2,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_20_20[7:0][7:0] = '{'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_20_21[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd2,3'd4},
'{3'd4,3'd2,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd2,3'd2,3'd4,3'd4,3'd2,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_20_22[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_20_23[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd3},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd3}};

parameter bit [2:0] SpriteTableR_20_24[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd1,3'd2,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd3,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd3,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_20_25[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd1,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd2,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd2,3'd1,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd3,3'd1,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd1,3'd4,3'd1},
'{3'd1,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_20_26[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd3,3'd2},
'{3'd4,3'd4,3'd1,3'd3,3'd2,3'd2,3'd3,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd1,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd1,3'd2,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd2,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4}};

parameter bit [2:0] SpriteTableR_20_27[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd3,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd1,3'd4}};

parameter bit [2:0] SpriteTableR_20_28[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd3,3'd4},
'{3'd3,3'd3,3'd1,3'd4,3'd1,3'd3,3'd1,3'd4},
'{3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd1,3'd4,3'd3,3'd2,3'd1,3'd1},
'{3'd4,3'd4,3'd1,3'd1,3'd4,3'd4,3'd2,3'd2},
'{3'd4,3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd2},
'{3'd3,3'd3,3'd1,3'd4,3'd3,3'd4,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_20_29[7:0][7:0] = '{'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd1,3'd4,3'd1},
'{3'd4,3'd3,3'd1,3'd4,3'd3,3'd3,3'd4,3'd3},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd1,3'd2,3'd1,3'd4,3'd1,3'd2,3'd1,3'd1},
'{3'd4,3'd1,3'd1,3'd1,3'd1,3'd3,3'd4,3'd4},
'{3'd4,3'd2,3'd1,3'd1,3'd1,3'd4,3'd3,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd3,3'd4,3'd3,3'd4}};

parameter bit [2:0] SpriteTableR_20_30[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd2,3'd4},
'{3'd1,3'd2,3'd1,3'd1,3'd1,3'd4,3'd2,3'd1},
'{3'd1,3'd2,3'd4,3'd1,3'd2,3'd1,3'd2,3'd1},
'{3'd1,3'd4,3'd2,3'd1,3'd3,3'd4,3'd3,3'd4},
'{3'd2,3'd4,3'd2,3'd4,3'd2,3'd4,3'd3,3'd3},
'{3'd4,3'd4,3'd2,3'd4,3'd2,3'd2,3'd1,3'd3},
'{3'd2,3'd4,3'd2,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd4,3'd2,3'd4,3'd2,3'd2,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_20_31[7:0][7:0] = '{'{3'd2,3'd4,3'd2,3'd4,3'd2,3'd2,3'd4,3'd4},
'{3'd2,3'd4,3'd2,3'd1,3'd4,3'd2,3'd4,3'd4},
'{3'd2,3'd4,3'd2,3'd4,3'd1,3'd2,3'd4,3'd2},
'{3'd2,3'd4,3'd1,3'd4,3'd4,3'd2,3'd4,3'd3},
'{3'd2,3'd4,3'd1,3'd4,3'd4,3'd2,3'd1,3'd3},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd2,3'd4,3'd1,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd2,3'd3,3'd4}};

parameter bit [2:0] SpriteTableR_20_32[7:0][7:0] = '{'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd4},
'{3'd3,3'd2,3'd4,3'd4,3'd4,3'd3,3'd3,3'd4},
'{3'd3,3'd3,3'd4,3'd4,3'd4,3'd3,3'd3,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd3,3'd2,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_20_33[7:0][7:0] = '{'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2},
'{3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_20_34[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd1}};

parameter bit [2:0] SpriteTableR_20_35[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd1,3'd1,3'd2,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_21_0[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_21_1[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_21_2[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_21_3[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_21_4[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2}};

parameter bit [2:0] SpriteTableR_21_5[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd1,3'd1},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd2,3'd4,3'd4,3'd4,3'd2}};

parameter bit [2:0] SpriteTableR_21_6[7:0][7:0] = '{'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd1,3'd2},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd1},
'{3'd3,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_21_7[7:0][7:0] = '{'{3'd3,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd3},
'{3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd2,3'd2,3'd2,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1}};

parameter bit [2:0] SpriteTableR_21_8[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd2,3'd1,3'd1,3'd2,3'd1,3'd1,3'd2,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd2,3'd1,3'd1,3'd2,3'd1,3'd1,3'd2,3'd1}};

parameter bit [2:0] SpriteTableR_21_9[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd2,3'd1,3'd1,3'd2,3'd1,3'd1,3'd2,3'd1},
'{3'd2,3'd1,3'd1,3'd2,3'd1,3'd1,3'd2,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd4,3'd1,3'd1,3'd4,3'd1,3'd1,3'd4,3'd1},
'{3'd2,3'd1,3'd1,3'd2,3'd1,3'd1,3'd2,3'd4},
'{3'd4,3'd1,3'd1,3'd4,3'd1,3'd1,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_21_10[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4},
'{3'd1,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd1,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4},
'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_21_11[7:0][7:0] = '{'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd2},
'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4},
'{3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2},
'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_21_12[7:0][7:0] = '{'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4},
'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4}};

parameter bit [2:0] SpriteTableR_21_13[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4},
'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd4,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2},
'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4}};

parameter bit [2:0] SpriteTableR_21_14[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4},
'{3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd4},
'{3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd4,3'd2,3'd4},
'{3'd2,3'd4,3'd4,3'd2,3'd1,3'd1,3'd2,3'd4},
'{3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_21_15[7:0][7:0] = '{'{3'd2,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd2,3'd2},
'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_21_16[7:0][7:0] = '{'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd2},
'{3'd2,3'd4,3'd4,3'd2,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd2,3'd4},
'{3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4},
'{3'd1,3'd1,3'd1,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_21_17[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd3},
'{3'd3,3'd3,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd1,3'd1,3'd1,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_21_18[7:0][7:0] = '{'{3'd1,3'd4,3'd4,3'd2,3'd4,3'd1,3'd1,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd1,3'd1,3'd4,3'd2,3'd1,3'd1,3'd2,3'd4},
'{3'd4,3'd1,3'd1,3'd1,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd1,3'd2,3'd4,3'd2,3'd2,3'd2},
'{3'd2,3'd4,3'd1,3'd2,3'd2,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_21_19[7:0][7:0] = '{'{3'd4,3'd1,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd2,3'd2,3'd4,3'd4},
'{3'd1,3'd1,3'd4,3'd2,3'd2,3'd3,3'd1,3'd1},
'{3'd1,3'd4,3'd4,3'd2,3'd4,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd2,3'd4,3'd1,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd2,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd2,3'd2,3'd4,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_21_20[7:0][7:0] = '{'{3'd2,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd2,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd2,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd2,3'd4,3'd4,3'd4,3'd3,3'd4},
'{3'd2,3'd2,3'd2,3'd4,3'd4,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_21_21[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2},
'{3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd4,3'd4,3'd2,3'd2,3'd4,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd1,3'd4,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_21_22[7:0][7:0] = '{'{3'd2,3'd2,3'd1,3'd4,3'd1,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd3,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_21_23[7:0][7:0] = '{'{3'd3,3'd1,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd1,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd3,3'd4,3'd2,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd1,3'd4,3'd3,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd1,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd3,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_21_24[7:0][7:0] = '{'{3'd1,3'd4,3'd4,3'd3,3'd4,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd1,3'd3,3'd4,3'd2,3'd2},
'{3'd4,3'd1,3'd4,3'd1,3'd4,3'd4,3'd2,3'd1},
'{3'd4,3'd3,3'd1,3'd4,3'd1,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd2},
'{3'd1,3'd2,3'd4,3'd4,3'd4,3'd3,3'd4,3'd2}};

parameter bit [2:0] SpriteTableR_21_25[7:0][7:0] = '{'{3'd1,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd1},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd1,3'd3,3'd4},
'{3'd3,3'd4,3'd4,3'd3,3'd4,3'd1,3'd1,3'd4},
'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd3}};

parameter bit [2:0] SpriteTableR_21_26[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd3,3'd4,3'd4},
'{3'd2,3'd2,3'd3,3'd1,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd2,3'd3,3'd4,3'd4,3'd3,3'd3,3'd1},
'{3'd3,3'd4,3'd4,3'd2,3'd1,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd2,3'd1,3'd4,3'd4,3'd2}};

parameter bit [2:0] SpriteTableR_21_27[7:0][7:0] = '{'{3'd4,3'd1,3'd2,3'd1,3'd1,3'd1,3'd2,3'd2},
'{3'd4,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2},
'{3'd1,3'd4,3'd4,3'd1,3'd1,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd2,3'd1,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd1,3'd1,3'd4,3'd4,3'd2},
'{3'd4,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd1,3'd1,3'd4,3'd2},
'{3'd1,3'd4,3'd2,3'd1,3'd1,3'd2,3'd4,3'd2}};

parameter bit [2:0] SpriteTableR_21_28[7:0][7:0] = '{'{3'd2,3'd4,3'd4,3'd1,3'd1,3'd4,3'd4,3'd2},
'{3'd3,3'd4,3'd4,3'd1,3'd1,3'd4,3'd4,3'd2},
'{3'd1,3'd2,3'd2,3'd2,3'd1,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd4,3'd4,3'd2,3'd2,3'd4,3'd4,3'd2},
'{3'd2,3'd4,3'd4,3'd2,3'd2,3'd4,3'd4,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_21_29[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd3,3'd4,3'd1},
'{3'd3,3'd4,3'd2,3'd4,3'd4,3'd3,3'd4,3'd1},
'{3'd3,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd1,3'd4,3'd4,3'd1,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_21_30[7:0][7:0] = '{'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd1,3'd3,3'd4},
'{3'd4,3'd3,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_21_31[7:0][7:0] = '{'{3'd1,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd2,3'd3,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd3,3'd2,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd2,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_21_32[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_21_33[7:0][7:0] = '{'{3'd1,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd1,3'd1,3'd4,3'd4},
'{3'd1,3'd2,3'd1,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd1,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1}};

parameter bit [2:0] SpriteTableR_21_34[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd1,3'd4,3'd2,3'd2,3'd2,3'd2,3'd1,3'd4}};

parameter bit [2:0] SpriteTableR_21_35[7:0][7:0] = '{'{3'd4,3'd1,3'd4,3'd2,3'd2,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd2,3'd2,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_22_0[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_22_1[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_22_2[7:0][7:0] = '{'{3'd4,3'd4,3'd2,3'd1,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd2,3'd2,3'd1,3'd1,3'd2,3'd2},
'{3'd1,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd1},
'{3'd1,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd1},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1},
'{3'd1,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_22_3[7:0][7:0] = '{'{3'd4,3'd1,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1},
'{3'd4,3'd1,3'd2,3'd1,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_22_4[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd1,3'd3},
'{3'd4,3'd1,3'd1,3'd1,3'd4,3'd4,3'd1,3'd4},
'{3'd1,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd1,3'd4,3'd4,3'd4,3'd1},
'{3'd2,3'd2,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd3,3'd4,3'd4,3'd4,3'd2}};

parameter bit [2:0] SpriteTableR_22_5[7:0][7:0] = '{'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd1,3'd1,3'd4,3'd4,3'd4,3'd1},
'{3'd2,3'd2,3'd4,3'd4,3'd1,3'd4,3'd3,3'd4},
'{3'd4,3'd2,3'd4,3'd4,3'd1,3'd4,3'd2,3'd4},
'{3'd4,3'd1,3'd2,3'd4,3'd4,3'd4,3'd1,3'd3},
'{3'd1,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd1,3'd4,3'd1,3'd4}};

parameter bit [2:0] SpriteTableR_22_6[7:0][7:0] = '{'{3'd2,3'd2,3'd4,3'd4,3'd2,3'd2,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd2,3'd2,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd2,3'd2,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd1,3'd4,3'd4,3'd4,3'd2,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd1,3'd4,3'd2,3'd3}};

parameter bit [2:0] SpriteTableR_22_7[7:0][7:0] = '{'{3'd4,3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd3,3'd2,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd2,3'd2,3'd1,3'd1,3'd2,3'd2},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd4,3'd3},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd4,3'd3}};

parameter bit [2:0] SpriteTableR_22_8[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd4,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd4,3'd4},
'{3'd1,3'd2,3'd1,3'd1,3'd1,3'd2,3'd2,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd4,3'd3,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd4,3'd3,3'd4},
'{3'd1,3'd2,3'd1,3'd1,3'd2,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_22_9[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd1,3'd2,3'd4,3'd4,3'd1,3'd4,3'd1,3'd4},
'{3'd1,3'd2,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd4,3'd4,3'd2,3'd2,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd2,3'd3,3'd4,3'd4},
'{3'd1,3'd2,3'd2,3'd1,3'd4,3'd3,3'd4,3'd4},
'{3'd1,3'd4,3'd1,3'd1,3'd4,3'd3,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_22_10[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd2,3'd1,3'd2,3'd4,3'd1,3'd4,3'd4},
'{3'd1,3'd4,3'd1,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd2,3'd3,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_22_11[7:0][7:0] = '{'{3'd4,3'd2,3'd2,3'd4,3'd3,3'd4,3'd4,3'd1},
'{3'd4,3'd2,3'd2,3'd4,3'd3,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd2,3'd1,3'd1,3'd4,3'd3}};

parameter bit [2:0] SpriteTableR_22_12[7:0][7:0] = '{'{3'd4,3'd2,3'd4,3'd3,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd3,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4},
'{3'd4,3'd2,3'd4,3'd1,3'd4,3'd4,3'd3,3'd4},
'{3'd4,3'd2,3'd4,3'd1,3'd4,3'd4,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_22_13[7:0][7:0] = '{'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd2,3'd4,3'd4,3'd1,3'd1,3'd4,3'd2},
'{3'd4,3'd4,3'd2,3'd4,3'd1,3'd4,3'd4,3'd2},
'{3'd4,3'd2,3'd2,3'd4,3'd4,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd3,3'd4,3'd2},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd3,3'd4,3'd1,3'd4,3'd2,3'd2},
'{3'd4,3'd4,3'd3,3'd4,3'd1,3'd4,3'd2,3'd4}};

parameter bit [2:0] SpriteTableR_22_14[7:0][7:0] = '{'{3'd4,3'd4,3'd3,3'd4,3'd3,3'd4,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd2,3'd2},
'{3'd4,3'd4,3'd1,3'd4,3'd3,3'd4,3'd4,3'd2},
'{3'd2,3'd4,3'd1,3'd4,3'd2,3'd2,3'd4,3'd2},
'{3'd2,3'd4,3'd4,3'd1,3'd4,3'd2,3'd4,3'd2},
'{3'd2,3'd4,3'd1,3'd1,3'd4,3'd2,3'd4,3'd2},
'{3'd2,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd2},
'{3'd2,3'd4,3'd1,3'd3,3'd4,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_22_15[7:0][7:0] = '{'{3'd2,3'd4,3'd1,3'd1,3'd1,3'd2,3'd2,3'd2},
'{3'd2,3'd3,3'd4,3'd4,3'd1,3'd4,3'd4,3'd2},
'{3'd4,3'd3,3'd1,3'd1,3'd1,3'd4,3'd4,3'd2},
'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd1,3'd2,3'd2},
'{3'd4,3'd3,3'd4,3'd3,3'd4,3'd1,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd3,3'd2,3'd3,3'd4,3'd1,3'd2,3'd2},
'{3'd4,3'd3,3'd2,3'd2,3'd4,3'd4,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_22_16[7:0][7:0] = '{'{3'd4,3'd1,3'd2,3'd2,3'd4,3'd1,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd2,3'd2,3'd2,3'd4,3'd2},
'{3'd1,3'd3,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd3,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd3,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd4,3'd2,3'd4,3'd3,3'd4,3'd3},
'{3'd4,3'd1,3'd1,3'd4,3'd1,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_22_17[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd1,3'd1,3'd1,3'd1,3'd4,3'd4},
'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_22_18[7:0][7:0] = '{'{3'd1,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd4,3'd4,3'd2,3'd1,3'd4,3'd2},
'{3'd4,3'd1,3'd1,3'd1,3'd1,3'd1,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_22_19[7:0][7:0] = '{'{3'd4,3'd1,3'd4,3'd4,3'd3,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd3},
'{3'd4,3'd3,3'd3,3'd3,3'd1,3'd1,3'd4,3'd3},
'{3'd2,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd3,3'd4,3'd1,3'd4,3'd3,3'd4},
'{3'd4,3'd3,3'd4,3'd4,3'd1,3'd1,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_22_20[7:0][7:0] = '{'{3'd4,3'd1,3'd4,3'd1,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd2,3'd4,3'd2},
'{3'd4,3'd3,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2},
'{3'd3,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2},
'{3'd2,3'd2,3'd2,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2}};

parameter bit [2:0] SpriteTableR_22_21[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd4,3'd1,3'd4},
'{3'd2,3'd2,3'd2,3'd4,3'd2,3'd1,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_22_22[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd1,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd3,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_22_23[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_22_24[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd4,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd1,3'd4,3'd1,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd1,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_22_25[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd2,3'd1,3'd2,3'd4,3'd3,3'd4,3'd1},
'{3'd4,3'd2,3'd1,3'd4,3'd1,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_22_26[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4},
'{3'd4,3'd4,3'd1,3'd3,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd2,3'd2,3'd4,3'd4},
'{3'd4,3'd3,3'd4,3'd4,3'd2,3'd4,3'd2,3'd4}};

parameter bit [2:0] SpriteTableR_22_27[7:0][7:0] = '{'{3'd2,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd2,3'd2,3'd2,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd4,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_22_28[7:0][7:0] = '{'{3'd2,3'd2,3'd4,3'd4,3'd2,3'd4,3'd2,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd2,3'd4,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd2,3'd2},
'{3'd2,3'd2,3'd4,3'd4,3'd2,3'd4,3'd2,3'd4},
'{3'd2,3'd2,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_22_29[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4},
'{3'd2,3'd1,3'd2,3'd2,3'd4,3'd2,3'd4,3'd4},
'{3'd2,3'd1,3'd2,3'd2,3'd4,3'd4,3'd2,3'd1},
'{3'd2,3'd1,3'd2,3'd2,3'd4,3'd4,3'd2,3'd3},
'{3'd4,3'd1,3'd1,3'd1,3'd4,3'd2,3'd4,3'd3},
'{3'd4,3'd1,3'd1,3'd1,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd1,3'd4,3'd2,3'd1,3'd3,3'd1},
'{3'd4,3'd4,3'd1,3'd2,3'd4,3'd1,3'd3,3'd4}};

parameter bit [2:0] SpriteTableR_22_30[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd2,3'd1,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd2,3'd1,3'd3,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd3,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd1}};

parameter bit [2:0] SpriteTableR_22_31[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2},
'{3'd4,3'd4,3'd1,3'd1,3'd1,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_22_32[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd1,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_22_33[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_22_34[7:0][7:0] = '{'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_22_35[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_23_0[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_23_1[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_23_2[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd1,3'd4,3'd4,3'd1,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_23_3[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_23_4[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd1,3'd2,3'd3,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd3,3'd3,3'd4,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_23_5[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd1,3'd4,3'd2,3'd1,3'd1,3'd2},
'{3'd3,3'd4,3'd1,3'd4,3'd4,3'd1,3'd1,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_23_6[7:0][7:0] = '{'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd2},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd1,3'd2,3'd3,3'd4,3'd4,3'd4},
'{3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd2,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd1,3'd4,3'd3}};

parameter bit [2:0] SpriteTableR_23_7[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd3,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd1,3'd1,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd3,3'd3,3'd2}};

parameter bit [2:0] SpriteTableR_23_8[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd2,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd1,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd2,3'd1,3'd1}};

parameter bit [2:0] SpriteTableR_23_9[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd1,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd1,3'd1,3'd1},
'{3'd4,3'd4,3'd1,3'd4,3'd2,3'd2,3'd1,3'd1},
'{3'd4,3'd4,3'd3,3'd4,3'd1,3'd2,3'd1,3'd1},
'{3'd4,3'd4,3'd3,3'd4,3'd1,3'd1,3'd1,3'd1},
'{3'd4,3'd4,3'd3,3'd4,3'd1,3'd1,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd2,3'd1,3'd2,3'd2,3'd1},
'{3'd4,3'd4,3'd4,3'd2,3'd1,3'd4,3'd1,3'd1}};

parameter bit [2:0] SpriteTableR_23_10[7:0][7:0] = '{'{3'd4,3'd1,3'd4,3'd2,3'd1,3'd1,3'd1,3'd1},
'{3'd4,3'd1,3'd4,3'd2,3'd1,3'd2,3'd4,3'd1},
'{3'd4,3'd3,3'd4,3'd4,3'd1,3'd2,3'd4,3'd1},
'{3'd4,3'd3,3'd4,3'd1,3'd1,3'd4,3'd1,3'd4},
'{3'd4,3'd2,3'd4,3'd1,3'd4,3'd2,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd4},
'{3'd1,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_23_11[7:0][7:0] = '{'{3'd3,3'd4,3'd2,3'd4,3'd4,3'd2,3'd2,3'd4},
'{3'd3,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd3,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4},
'{3'd4,3'd2,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4},
'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4}};

parameter bit [2:0] SpriteTableR_23_12[7:0][7:0] = '{'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd1,3'd2,3'd2},
'{3'd4,3'd4,3'd2,3'd2,3'd4,3'd1,3'd2,3'd4}};

parameter bit [2:0] SpriteTableR_23_13[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4},
'{3'd2,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_23_14[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_23_15[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_23_16[7:0][7:0] = '{'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd3,3'd3,3'd4,3'd1,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2}};

parameter bit [2:0] SpriteTableR_23_17[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd3,3'd3,3'd3,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd2,3'd2,3'd4,3'd2,3'd1},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd1,3'd1,3'd4,3'd4,3'd2},
'{3'd1,3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_23_18[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd2,3'd1,3'd4,3'd2,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_23_19[7:0][7:0] = '{'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4},
'{3'd4,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2}};

parameter bit [2:0] SpriteTableR_23_20[7:0][7:0] = '{'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4},
'{3'd4,3'd4,3'd2,3'd2,3'd4,3'd2,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd1},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd4,3'd3,3'd4},
'{3'd2,3'd4,3'd2,3'd2,3'd2,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4},
'{3'd2,3'd4,3'd2,3'd4,3'd3,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_23_21[7:0][7:0] = '{'{3'd2,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd1,3'd1,3'd4,3'd4,3'd1,3'd4},
'{3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd3,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_23_22[7:0][7:0] = '{'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_23_23[7:0][7:0] = '{'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd2},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd3,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd1,3'd1,3'd1,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd3,3'd4,3'd4,3'd3,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_23_24[7:0][7:0] = '{'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd2,3'd2,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4},
'{3'd2,3'd2,3'd2,3'd4,3'd1,3'd1,3'd4,3'd3},
'{3'd2,3'd2,3'd2,3'd4,3'd3,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd3,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_23_25[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd2,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd1,3'd4},
'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_23_26[7:0][7:0] = '{'{3'd3,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3},
'{3'd4,3'd4,3'd4,3'd2,3'd1,3'd1,3'd4,3'd4},
'{3'd4,3'd2,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd1,3'd4,3'd4,3'd1,3'd4,3'd3},
'{3'd4,3'd1,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd1,3'd4,3'd2,3'd1,3'd4,3'd3}};

parameter bit [2:0] SpriteTableR_23_27[7:0][7:0] = '{'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd3,3'd3,3'd4,3'd4,3'd1},
'{3'd2,3'd4,3'd1,3'd4,3'd4,3'd1,3'd4,3'd3},
'{3'd2,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_23_28[7:0][7:0] = '{'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd2,3'd4,3'd4,3'd2,3'd2,3'd1,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd2,3'd4,3'd4,3'd2,3'd2,3'd2,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd2,3'd2,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd1,3'd4,3'd1,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_23_29[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_23_30[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_23_31[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd1,3'd4,3'd4,3'd1,3'd1,3'd1},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd1,3'd4},
'{3'd2,3'd4,3'd4,3'd2,3'd2,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd2,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd2,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_23_32[7:0][7:0] = '{'{3'd1,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd2,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd2,3'd1,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd1,3'd1,3'd2,3'd1,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd1,3'd1,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_23_33[7:0][7:0] = '{'{3'd1,3'd4,3'd4,3'd2,3'd1,3'd1,3'd2,3'd2},
'{3'd2,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd2,3'd2,3'd2,3'd4},
'{3'd4,3'd2,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_23_34[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd1,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd2,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_23_35[7:0][7:0] = '{'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1},
'{3'd4,3'd1,3'd2,3'd2,3'd2,3'd2,3'd1,3'd4},
'{3'd4,3'd1,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_24_0[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd1,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_24_1[7:0][7:0] = '{'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_24_2[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd4,3'd4,3'd2,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd1,3'd4,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_24_3[7:0][7:0] = '{'{3'd2,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_24_4[7:0][7:0] = '{'{3'd4,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd3,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1},
'{3'd1,3'd4,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd2,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd2,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd1,3'd4,3'd3,3'd3,3'd4,3'd4},
'{3'd2,3'd1,3'd4,3'd4,3'd3,3'd3,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_24_5[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd2,3'd2,3'd3,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd2,3'd4,3'd2,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd1,3'd2,3'd1,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_24_6[7:0][7:0] = '{'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd3,3'd4,3'd1,3'd4,3'd4,3'd1,3'd4},
'{3'd2,3'd1,3'd4,3'd4,3'd3,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd4},
'{3'd4,3'd3,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd3,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd2,3'd1,3'd4}};

parameter bit [2:0] SpriteTableR_24_7[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd1,3'd1,3'd4,3'd3,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_24_8[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd2,3'd1,3'd1,3'd2,3'd1,3'd1,3'd2,3'd1}};

parameter bit [2:0] SpriteTableR_24_9[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd2,3'd1,3'd1,3'd2,3'd1,3'd1,3'd2,3'd1},
'{3'd2,3'd1,3'd1,3'd2,3'd1,3'd1,3'd2,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2},
'{3'd2,3'd2,3'd1,3'd2,3'd2,3'd1,3'd2,3'd2},
'{3'd1,3'd1,3'd1,3'd1,3'd4,3'd1,3'd1,3'd2}};

parameter bit [2:0] SpriteTableR_24_10[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd2,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1,3'd4},
'{3'd2,3'd2,3'd1,3'd2,3'd1,3'd1,3'd1,3'd4},
'{3'd4,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd4},
'{3'd2,3'd1,3'd1,3'd1,3'd4,3'd1,3'd1,3'd3},
'{3'd2,3'd2,3'd1,3'd1,3'd2,3'd1,3'd2,3'd3},
'{3'd4,3'd1,3'd1,3'd1,3'd4,3'd1,3'd2,3'd3},
'{3'd4,3'd1,3'd1,3'd1,3'd4,3'd4,3'd4,3'd3}};

parameter bit [2:0] SpriteTableR_24_11[7:0][7:0] = '{'{3'd2,3'd2,3'd1,3'd1,3'd2,3'd1,3'd4,3'd3},
'{3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1},
'{3'd4,3'd1,3'd1,3'd1,3'd4,3'd2,3'd2,3'd3},
'{3'd2,3'd2,3'd1,3'd2,3'd4,3'd2,3'd4,3'd2},
'{3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd1,3'd1,3'd1,3'd1,3'd4},
'{3'd2,3'd2,3'd1,3'd2,3'd2,3'd1,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_24_12[7:0][7:0] = '{'{3'd2,3'd2,3'd1,3'd2,3'd2,3'd4,3'd2,3'd2},
'{3'd4,3'd4,3'd1,3'd1,3'd4,3'd1,3'd1,3'd4},
'{3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2},
'{3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd2,3'd4,3'd2,3'd3,3'd3},
'{3'd2,3'd2,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_24_13[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd2,3'd4,3'd1,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd2,3'd4,3'd4,3'd4,3'd1},
'{3'd2,3'd4,3'd4,3'd2,3'd2,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd3,3'd4,3'd4,3'd3},
'{3'd2,3'd2,3'd4,3'd4,3'd3,3'd4,3'd4,3'd3},
'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd2,3'd4,3'd2,3'd4,3'd1,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_24_14[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd4,3'd1,3'd4,3'd1,3'd4},
'{3'd2,3'd2,3'd2,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd2,3'd3,3'd4,3'd4,3'd4,3'd3},
'{3'd2,3'd2,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd3,3'd1,3'd4,3'd4,3'd1},
'{3'd2,3'd2,3'd4,3'd1,3'd4,3'd4,3'd4,3'd1},
'{3'd2,3'd2,3'd4,3'd4,3'd3,3'd3,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2}};

parameter bit [2:0] SpriteTableR_24_15[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd1,3'd1},
'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2},
'{3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_24_16[7:0][7:0] = '{'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2},
'{3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd3},
'{3'd3,3'd3,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd1,3'd4,3'd3,3'd3,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_24_17[7:0][7:0] = '{'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd3,3'd4,3'd4,3'd3,3'd3,3'd4,3'd1},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_24_18[7:0][7:0] = '{'{3'd2,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd3,3'd4,3'd4},
'{3'd2,3'd4,3'd3,3'd4,3'd4,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd3,3'd4,3'd4},
'{3'd4,3'd2,3'd3,3'd4,3'd4,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd3,3'd4,3'd4},
'{3'd2,3'd4,3'd3,3'd4,3'd4,3'd3,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_24_19[7:0][7:0] = '{'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd3,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd2,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_24_20[7:0][7:0] = '{'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_24_21[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd3,3'd1},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd3,3'd1,3'd1,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_24_22[7:0][7:0] = '{'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_24_23[7:0][7:0] = '{'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd2,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd1,3'd2,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_24_24[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd3,3'd4,3'd1,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_24_25[7:0][7:0] = '{'{3'd4,3'd4,3'd2,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd2,3'd2,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd1,3'd2,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd3,3'd1,3'd1},
'{3'd3,3'd1,3'd3,3'd4,3'd4,3'd4,3'd2,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4}};

parameter bit [2:0] SpriteTableR_24_26[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd3,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd2,3'd3,3'd4,3'd4},
'{3'd4,3'd3,3'd4,3'd1,3'd4,3'd4,3'd1,3'd4},
'{3'd2,3'd1,3'd4,3'd4,3'd3,3'd3,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_24_27[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd1,3'd4,3'd4,3'd1,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4}};

parameter bit [2:0] SpriteTableR_24_28[7:0][7:0] = '{'{3'd4,3'd1,3'd4,3'd4,3'd2,3'd2,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd1,3'd2,3'd2,3'd1,3'd1},
'{3'd1,3'd3,3'd3,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_24_29[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_24_30[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_24_31[7:0][7:0] = '{'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_24_32[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd1,3'd1,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_24_33[7:0][7:0] = '{'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1},
'{3'd4,3'd2,3'd3,3'd1,3'd4,3'd1,3'd2,3'd4},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd4,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd1},
'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd1,3'd1},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4}};

parameter bit [2:0] SpriteTableR_24_34[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_24_35[7:0][7:0] = '{'{3'd1,3'd4,3'd4,3'd1,3'd4,3'd4,3'd1,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_25_0[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_25_1[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd1,3'd1},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_25_2[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd2,3'd1},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_25_3[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd1,3'd4,3'd1,3'd1,3'd2,3'd2,3'd2},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4}};

parameter bit [2:0] SpriteTableR_25_4[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd3,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4}};

parameter bit [2:0] SpriteTableR_25_5[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd1,3'd2,3'd1,3'd4,3'd4,3'd1,3'd2,3'd1},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd2,3'd2,3'd1},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_25_6[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd4},
'{3'd3,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd3,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd1,3'd4,3'd4,3'd2,3'd1,3'd4},
'{3'd2,3'd4,3'd2,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_25_7[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd4},
'{3'd3,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1}};

parameter bit [2:0] SpriteTableR_25_8[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1}};

parameter bit [2:0] SpriteTableR_25_9[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_25_10[7:0][7:0] = '{'{3'd3,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd3,3'd4,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd2,3'd4},
'{3'd1,3'd4,3'd4,3'd3,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd1,3'd2,3'd2,3'd3,3'd3,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_25_11[7:0][7:0] = '{'{3'd4,3'd1,3'd1,3'd4,3'd1,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd1},
'{3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd2,3'd3},
'{3'd2,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2},
'{3'd4,3'd1,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd1,3'd4,3'd1,3'd1,3'd1},
'{3'd4,3'd2,3'd2,3'd1,3'd2,3'd2,3'd1,3'd2}};

parameter bit [2:0] SpriteTableR_25_12[7:0][7:0] = '{'{3'd4,3'd2,3'd2,3'd1,3'd2,3'd2,3'd1,3'd1},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd4},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2},
'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd3,3'd4,3'd3,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_25_13[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd1,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_25_14[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd1,3'd4,3'd1,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd4,3'd4},
'{3'd4,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd4,3'd1},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_25_15[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd1},
'{3'd4,3'd2,3'd2,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd2,3'd2,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd3,3'd1},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd4,3'd3,3'd4},
'{3'd4,3'd2,3'd2,3'd4,3'd4,3'd4,3'd3,3'd4},
'{3'd2,3'd2,3'd2,3'd4,3'd2,3'd4,3'd3,3'd4},
'{3'd4,3'd2,3'd2,3'd4,3'd2,3'd4,3'd3,3'd4}};

parameter bit [2:0] SpriteTableR_25_16[7:0][7:0] = '{'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd3,3'd3,3'd4,3'd1,3'd4},
'{3'd1,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd3,3'd2},
'{3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3}};

parameter bit [2:0] SpriteTableR_25_17[7:0][7:0] = '{'{3'd4,3'd1,3'd3,3'd4,3'd1,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4}};

parameter bit [2:0] SpriteTableR_25_18[7:0][7:0] = '{'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd1,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd2,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_25_19[7:0][7:0] = '{'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_25_20[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd1,3'd4,3'd1,3'd1,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_25_21[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd1,3'd3,3'd4,3'd2,3'd2,3'd2},
'{3'd1,3'd3,3'd3,3'd1,3'd4,3'd1,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_25_22[7:0][7:0] = '{'{3'd4,3'd1,3'd3,3'd3,3'd1,3'd1,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd3,3'd3,3'd4,3'd1,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd1,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd2,3'd3,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd3,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_25_23[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd3,3'd3,3'd4},
'{3'd4,3'd3,3'd4,3'd3,3'd1,3'd4,3'd3,3'd3},
'{3'd1,3'd4,3'd4,3'd1,3'd3,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd3,3'd4,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd2,3'd4,3'd4,3'd3},
'{3'd4,3'd2,3'd2,3'd4,3'd4,3'd2,3'd2,3'd2},
'{3'd4,3'd2,3'd4,3'd2,3'd2,3'd2,3'd4,3'd2}};

parameter bit [2:0] SpriteTableR_25_24[7:0][7:0] = '{'{3'd1,3'd4,3'd2,3'd2,3'd2,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd2,3'd2,3'd4,3'd4,3'd2},
'{3'd4,3'd1,3'd4,3'd2,3'd2,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd2,3'd2,3'd4,3'd2,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_25_25[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd2,3'd2,3'd2,3'd2,3'd1,3'd4,3'd4},
'{3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4},
'{3'd4,3'd2,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_25_26[7:0][7:0] = '{'{3'd2,3'd4,3'd2,3'd1,3'd4,3'd3,3'd3,3'd4},
'{3'd3,3'd4,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd2,3'd4,3'd4,3'd1,3'd1,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd3,3'd1,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd3},
'{3'd1,3'd4,3'd4,3'd4,3'd3,3'd2,3'd3,3'd4}};

parameter bit [2:0] SpriteTableR_25_27[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd3,3'd3,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_25_28[7:0][7:0] = '{'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd1,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3}};

parameter bit [2:0] SpriteTableR_25_29[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_25_30[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_25_31[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_25_32[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_25_33[7:0][7:0] = '{'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd4,3'd4,3'd1,3'd3},
'{3'd4,3'd4,3'd1,3'd1,3'd1,3'd2,3'd2,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_25_34[7:0][7:0] = '{'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_25_35[7:0][7:0] = '{'{3'd2,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_26_0[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_26_1[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_26_2[7:0][7:0] = '{'{3'd4,3'd1,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_26_3[7:0][7:0] = '{'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_26_4[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_26_5[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd3,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd4,3'd4,3'd4,3'd1,3'd1},
'{3'd1,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_26_6[7:0][7:0] = '{'{3'd4,3'd1,3'd2,3'd4,3'd4,3'd4,3'd1,3'd1},
'{3'd4,3'd1,3'd4,3'd1,3'd4,3'd4,3'd1,3'd1},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1}};

parameter bit [2:0] SpriteTableR_26_7[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1},
'{3'd3,3'd3,3'd3,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd2,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd4}};

parameter bit [2:0] SpriteTableR_26_8[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd4,3'd3},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd4,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd4}};

parameter bit [2:0] SpriteTableR_26_9[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd2,3'd1,3'd4,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_26_10[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd3,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd2,3'd1,3'd4,3'd2,3'd2},
'{3'd2,3'd4,3'd2,3'd2,3'd2,3'd2,3'd1,3'd4},
'{3'd1,3'd4,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_26_11[7:0][7:0] = '{'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd4,3'd4,3'd3,3'd4,3'd2},
'{3'd3,3'd4,3'd3,3'd4,3'd4,3'd4,3'd2,3'd2},
'{3'd2,3'd4,3'd3,3'd4,3'd4,3'd3,3'd4,3'd4},
'{3'd2,3'd4,3'd3,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd1,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd1,3'd1,3'd1,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_26_12[7:0][7:0] = '{'{3'd2,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd3,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_26_13[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_26_14[7:0][7:0] = '{'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_26_15[7:0][7:0] = '{'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd2,3'd3},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_26_16[7:0][7:0] = '{'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd3,3'd4,3'd4},
'{3'd3,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_26_17[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_26_18[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd1,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_26_19[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_26_20[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd3,3'd3,3'd3,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_26_21[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd1,3'd2}};

parameter bit [2:0] SpriteTableR_26_22[7:0][7:0] = '{'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd1,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd2,3'd2},
'{3'd3,3'd3,3'd4,3'd1,3'd2,3'd1,3'd4,3'd4},
'{3'd3,3'd3,3'd3,3'd1,3'd4,3'd3,3'd2,3'd1},
'{3'd1,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_26_23[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd2,3'd3,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd2},
'{3'd3,3'd3,3'd4,3'd4,3'd4,3'd2,3'd2,3'd4},
'{3'd4,3'd3,3'd3,3'd4,3'd3,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd3,3'd3,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd3,3'd2,3'd4,3'd4,3'd4},
'{3'd2,3'd1,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_26_24[7:0][7:0] = '{'{3'd2,3'd2,3'd1,3'd2,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd1,3'd4,3'd4},
'{3'd2,3'd4,3'd2,3'd3,3'd3,3'd3,3'd4,3'd4},
'{3'd3,3'd1,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_26_25[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_26_26[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd4,3'd1,3'd1,3'd4,3'd3,3'd3},
'{3'd4,3'd1,3'd4,3'd4,3'd3,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd1,3'd1,3'd4,3'd4,3'd1,3'd4,3'd1,3'd2}};

parameter bit [2:0] SpriteTableR_26_27[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd1,3'd1},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_26_28[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd1,3'd3,3'd3,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_26_29[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_26_30[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_26_31[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_26_32[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd1,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_26_33[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd3,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_26_34[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_26_35[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_27_0[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_27_1[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_27_2[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_27_3[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd2},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd1,3'd4,3'd1,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd1,3'd1,3'd2},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_27_4[7:0][7:0] = '{'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_27_5[7:0][7:0] = '{'{3'd4,3'd4,3'd1,3'd2,3'd2,3'd2,3'd2,3'd1},
'{3'd4,3'd4,3'd1,3'd2,3'd2,3'd2,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd2,3'd2,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd2,3'd2,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd2,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4}};

parameter bit [2:0] SpriteTableR_27_6[7:0][7:0] = '{'{3'd1,3'd1,3'd4,3'd1,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd2,3'd2,3'd4,3'd1},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd1,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd4}};

parameter bit [2:0] SpriteTableR_27_7[7:0][7:0] = '{'{3'd4,3'd4,3'd2,3'd2,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd2},
'{3'd1,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_27_8[7:0][7:0] = '{'{3'd1,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd3,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_27_9[7:0][7:0] = '{'{3'd4,3'd3,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd2,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd4}};

parameter bit [2:0] SpriteTableR_27_10[7:0][7:0] = '{'{3'd2,3'd4,3'd2,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd4,3'd1,3'd2,3'd2,3'd2,3'd4,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd1,3'd2,3'd4,3'd4,3'd4},
'{3'd1,3'd3,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_27_11[7:0][7:0] = '{'{3'd2,3'd4,3'd4,3'd2,3'd4,3'd4,3'd3,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd3,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd3,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_27_12[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_27_13[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_27_14[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_27_15[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd1,3'd4},
'{3'd1,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_27_16[7:0][7:0] = '{'{3'd4,3'd4,3'd1,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd3,3'd2,3'd4},
'{3'd4,3'd4,3'd1,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_27_17[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd1,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_27_18[7:0][7:0] = '{'{3'd4,3'd4,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2}};

parameter bit [2:0] SpriteTableR_27_19[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_27_20[7:0][7:0] = '{'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd4,3'd4,3'd2,3'd2,3'd1,3'd4},
'{3'd3,3'd4,3'd3,3'd4,3'd3,3'd2,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4}};

parameter bit [2:0] SpriteTableR_27_21[7:0][7:0] = '{'{3'd1,3'd1,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd4},
'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_27_22[7:0][7:0] = '{'{3'd4,3'd1,3'd1,3'd2,3'd2,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd1,3'd4,3'd2,3'd4,3'd3,3'd1},
'{3'd1,3'd4,3'd2,3'd4,3'd4,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd2,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_27_23[7:0][7:0] = '{'{3'd3,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_27_24[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_27_25[7:0][7:0] = '{'{3'd4,3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd3,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd2,3'd3,3'd2,3'd3,3'd3,3'd3},
'{3'd1,3'd4,3'd1,3'd4,3'd4,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_27_26[7:0][7:0] = '{'{3'd2,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd1,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_27_27[7:0][7:0] = '{'{3'd3,3'd1,3'd1,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd3,3'd2,3'd1,3'd1,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd1,3'd1,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_27_28[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_27_29[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_27_30[7:0][7:0] = '{'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd1,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_27_31[7:0][7:0] = '{'{3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_27_32[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd3},
'{3'd4,3'd4,3'd1,3'd1,3'd4,3'd4,3'd3,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_27_33[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2}};

parameter bit [2:0] SpriteTableR_27_34[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_27_35[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_28_0[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_28_1[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3}};

parameter bit [2:0] SpriteTableR_28_2[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd1,3'd2,3'd4,3'd3,3'd3},
'{3'd4,3'd4,3'd1,3'd4,3'd3,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_28_3[7:0][7:0] = '{'{3'd2,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd2,3'd3,3'd3,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd2,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd3,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_28_4[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd3,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd1,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd1,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_28_5[7:0][7:0] = '{'{3'd4,3'd1,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_28_6[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_28_7[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd4,3'd2,3'd1,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd1,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_28_8[7:0][7:0] = '{'{3'd2,3'd4,3'd4,3'd4,3'd2,3'd1,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd1,3'd2,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_28_9[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4},
'{3'd1,3'd1,3'd1,3'd4,3'd4,3'd4,3'd1,3'd2},
'{3'd4,3'd1,3'd4,3'd1,3'd4,3'd1,3'd1,3'd2},
'{3'd4,3'd1,3'd1,3'd1,3'd4,3'd2,3'd2,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd1,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd4,3'd4},
'{3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd4,3'd1},
'{3'd4,3'd1,3'd1,3'd2,3'd4,3'd1,3'd4,3'd2}};

parameter bit [2:0] SpriteTableR_28_10[7:0][7:0] = '{'{3'd4,3'd2,3'd1,3'd2,3'd4,3'd3,3'd1,3'd1},
'{3'd2,3'd2,3'd1,3'd1,3'd2,3'd1,3'd4,3'd4},
'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd1,3'd2},
'{3'd4,3'd1,3'd1,3'd1,3'd2,3'd4,3'd3,3'd3},
'{3'd4,3'd2,3'd4,3'd4,3'd1,3'd3,3'd2,3'd2},
'{3'd4,3'd4,3'd3,3'd3,3'd3,3'd2,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd1,3'd3,3'd2,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_28_11[7:0][7:0] = '{'{3'd1,3'd4,3'd4,3'd3,3'd4,3'd2,3'd2,3'd2},
'{3'd4,3'd1,3'd3,3'd4,3'd4,3'd4,3'd2,3'd2},
'{3'd4,3'd2,3'd2,3'd2,3'd4,3'd4,3'd4,3'd2},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd3,3'd1,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_28_12[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_28_13[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_28_14[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd2,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd2,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_28_15[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_28_16[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd2,3'd1,3'd1,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd1,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_28_17[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd1},
'{3'd4,3'd4,3'd2,3'd2,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_28_18[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd2,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1},
'{3'd4,3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1}};

parameter bit [2:0] SpriteTableR_28_19[7:0][7:0] = '{'{3'd4,3'd2,3'd2,3'd1,3'd4,3'd2,3'd4,3'd4},
'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd2,3'd2,3'd2,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd2,3'd2,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd3,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_28_20[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd1,3'd1},
'{3'd4,3'd1,3'd4,3'd4,3'd1,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd1,3'd1,3'd2,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_28_21[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2},
'{3'd4,3'd1,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_28_22[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd3,3'd4,3'd2,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_28_23[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_28_24[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_28_25[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd3,3'd4,3'd1,3'd4,3'd4},
'{3'd3,3'd4,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_28_26[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_28_27[7:0][7:0] = '{'{3'd4,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_28_28[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_28_29[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd3,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd3,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd3,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_28_30[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd1,3'd3,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd1,3'd4,3'd1,3'd1,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd1,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_28_31[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_28_32[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd3,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_28_33[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd4,3'd2,3'd1,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_28_34[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd1,3'd1,3'd2,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_28_35[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_29_0[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_29_1[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd3,3'd3,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd3,3'd1,3'd1,3'd1},
'{3'd4,3'd4,3'd1,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd3,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_29_2[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd1,3'd1,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_29_3[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_29_4[7:0][7:0] = '{'{3'd1,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3},
'{3'd4,3'd3,3'd2,3'd4,3'd1,3'd1,3'd3,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd1,3'd4}};

parameter bit [2:0] SpriteTableR_29_5[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_29_6[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd1,3'd1,3'd1,3'd1,3'd4},
'{3'd4,3'd2,3'd2,3'd4,3'd1,3'd1,3'd4,3'd4},
'{3'd4,3'd2,3'd2,3'd4,3'd1,3'd1,3'd4,3'd4},
'{3'd4,3'd2,3'd2,3'd1,3'd2,3'd2,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_29_7[7:0][7:0] = '{'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4},
'{3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd4},
'{3'd1,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4},
'{3'd1,3'd4,3'd2,3'd1,3'd4,3'd1,3'd1,3'd1},
'{3'd4,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_29_8[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_29_9[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd2,3'd2,3'd4,3'd2,3'd1},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4},
'{3'd2,3'd2,3'd1,3'd2,3'd1,3'd1,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_29_10[7:0][7:0] = '{'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd1,3'd2,3'd4,3'd2,3'd4},
'{3'd1,3'd2,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd1,3'd4},
'{3'd1,3'd1,3'd2,3'd4,3'd4,3'd1,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_29_11[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd2,3'd4}};

parameter bit [2:0] SpriteTableR_29_12[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd1,3'd2,3'd2,3'd1,3'd2},
'{3'd4,3'd4,3'd1,3'd2,3'd2,3'd2,3'd1,3'd2},
'{3'd4,3'd4,3'd1,3'd4,3'd1,3'd4,3'd2,3'd1},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd1,3'd4,3'd1,3'd2,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_29_13[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd1,3'd4,3'd1,3'd2,3'd1,3'd4},
'{3'd2,3'd4,3'd1,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd2,3'd4,3'd4,3'd1,3'd3,3'd4,3'd4},
'{3'd3,3'd4,3'd1,3'd4,3'd1,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_29_14[7:0][7:0] = '{'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd3,3'd4,3'd4,3'd4,3'd3,3'd1,3'd4},
'{3'd3,3'd4,3'd1,3'd4,3'd1,3'd4,3'd1,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_29_15[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd1},
'{3'd4,3'd4,3'd1,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_29_16[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd1,3'd1,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_29_17[7:0][7:0] = '{'{3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd2,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd2,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_29_18[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_29_19[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_29_20[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd4,3'd4,3'd1,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd1,3'd1,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd1,3'd4},
'{3'd4,3'd4,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd4,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_29_21[7:0][7:0] = '{'{3'd4,3'd1,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd2,3'd1,3'd1,3'd2,3'd2,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd1,3'd4,3'd4},
'{3'd1,3'd1,3'd2,3'd4,3'd2,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_29_22[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd2,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4}};

parameter bit [2:0] SpriteTableR_29_23[7:0][7:0] = '{'{3'd4,3'd2,3'd1,3'd1,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd2,3'd2,3'd2,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_29_24[7:0][7:0] = '{'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4}};

parameter bit [2:0] SpriteTableR_29_25[7:0][7:0] = '{'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd2},
'{3'd1,3'd1,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd1,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd1,3'd4,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd1,3'd4,3'd2,3'd2,3'd2,3'd1,3'd2,3'd2},
'{3'd4,3'd4,3'd2,3'd2,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_29_26[7:0][7:0] = '{'{3'd1,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd2,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd1,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd2,3'd1,3'd4}};

parameter bit [2:0] SpriteTableR_29_27[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_29_28[7:0][7:0] = '{'{3'd2,3'd4,3'd1,3'd1,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd1,3'd1,3'd1,3'd1,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_29_29[7:0][7:0] = '{'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd4,3'd4,3'd1,3'd1,3'd4,3'd4},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd3,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_29_30[7:0][7:0] = '{'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_29_31[7:0][7:0] = '{'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd1,3'd1,3'd1,3'd4,3'd4,3'd4},
'{3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_29_32[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_29_33[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_29_34[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_29_35[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_30_0[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_30_1[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd1,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_30_2[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1}};

parameter bit [2:0] SpriteTableR_30_3[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd3},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd3},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd3,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd1,3'd3,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_30_4[7:0][7:0] = '{'{3'd4,3'd1,3'd4,3'd2,3'd1,3'd4,3'd4,3'd4},
'{3'd3,3'd2,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd1,3'd4,3'd4,3'd4},
'{3'd2,3'd1,3'd4,3'd1,3'd4,3'd1,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_30_5[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_30_6[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_30_7[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd2,3'd1,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd1,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd1,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_30_8[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd2,3'd1,3'd4},
'{3'd4,3'd4,3'd2,3'd2,3'd2,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd2,3'd2,3'd1,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd4,3'd1,3'd2,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_30_9[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_30_10[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_30_11[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd1},
'{3'd1,3'd1,3'd1,3'd4,3'd1,3'd2,3'd2,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd2,3'd1},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd4,3'd4,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableR_30_12[7:0][7:0] = '{'{3'd2,3'd1,3'd2,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd2,3'd2},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd2,3'd2,3'd2},
'{3'd4,3'd1,3'd1,3'd4,3'd4,3'd2,3'd2,3'd1},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_30_13[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_30_14[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd3,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd1,3'd1,3'd4,3'd1,3'd1,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_30_15[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1},
'{3'd4,3'd2,3'd2,3'd2,3'd4,3'd2,3'd1,3'd1},
'{3'd1,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_30_16[7:0][7:0] = '{'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_30_17[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd1,3'd1,3'd1,3'd4},
'{3'd4,3'd1,3'd2,3'd1,3'd1,3'd1,3'd4,3'd4},
'{3'd4,3'd1,3'd2,3'd2,3'd2,3'd1,3'd4,3'd4},
'{3'd1,3'd2,3'd2,3'd1,3'd4,3'd1,3'd4,3'd4},
'{3'd1,3'd2,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1}};

parameter bit [2:0] SpriteTableR_30_18[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_30_19[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd1,3'd1,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_30_20[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd2,3'd1,3'd1,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_30_21[7:0][7:0] = '{'{3'd4,3'd2,3'd2,3'd2,3'd1,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_30_22[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_30_23[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_30_24[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_30_25[7:0][7:0] = '{'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_30_26[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_30_27[7:0][7:0] = '{'{3'd4,3'd4,3'd1,3'd1,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_30_28[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_30_29[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_30_30[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_30_31[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_30_32[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_30_33[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_30_34[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_30_35[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_31_0[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_31_1[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd1,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_31_2[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd2,3'd1,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd3,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd3,3'd3,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd3,3'd3,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd3,3'd3,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd2,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_31_3[7:0][7:0] = '{'{3'd4,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd3,3'd3,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd3,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_31_4[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_31_5[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_31_6[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_31_7[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_31_8[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_31_9[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_31_10[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_31_11[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_31_12[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd1,3'd4,3'd1,3'd4,3'd4},
'{3'd2,3'd2,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd2,3'd4,3'd1,3'd4,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd4,3'd4},
'{3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd4},
'{3'd4,3'd4,3'd2,3'd1,3'd1,3'd1,3'd4,3'd4},
'{3'd4,3'd1,3'd2,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_31_13[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_31_14[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_31_15[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_31_16[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_31_17[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_31_18[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_31_19[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_31_20[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_31_21[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_31_22[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_31_23[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_31_24[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_31_25[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_31_26[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_31_27[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_31_28[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_31_29[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_31_30[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_31_31[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_31_32[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_31_33[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_31_34[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableR_31_35[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

logic [9:0] SpriteTableG;

parameter bit [7:0] SpritePaletteG[4:0] = '{8'd255, 8'd183, 8'd151, 8'd8, 8'd222};

	always_comb
	begin
		SpriteTableG = 10'd0;
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableG = SpriteTableG_0_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableG = SpriteTableG_0_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableG = SpriteTableG_0_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableG = SpriteTableG_0_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableG = SpriteTableG_0_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableG = SpriteTableG_0_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableG = SpriteTableG_0_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableG = SpriteTableG_0_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableG = SpriteTableG_0_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableG = SpriteTableG_0_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableG = SpriteTableG_0_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableG = SpriteTableG_0_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableG = SpriteTableG_0_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_0_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableG = SpriteTableG_0_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableG = SpriteTableG_0_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableG = SpriteTableG_0_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableG = SpriteTableG_0_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableG = SpriteTableG_0_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableG = SpriteTableG_0_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableG = SpriteTableG_0_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableG = SpriteTableG_0_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableG = SpriteTableG_0_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableG = SpriteTableG_0_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableG = SpriteTableG_0_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableG = SpriteTableG_0_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableG = SpriteTableG_0_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableG = SpriteTableG_0_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableG = SpriteTableG_0_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableG = SpriteTableG_0_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableG = SpriteTableG_0_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableG = SpriteTableG_0_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableG = SpriteTableG_0_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableG = SpriteTableG_0_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableG = SpriteTableG_0_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableG = SpriteTableG_0_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableG = SpriteTableG_1_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableG = SpriteTableG_1_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableG = SpriteTableG_1_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableG = SpriteTableG_1_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableG = SpriteTableG_1_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableG = SpriteTableG_1_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableG = SpriteTableG_1_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableG = SpriteTableG_1_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableG = SpriteTableG_1_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableG = SpriteTableG_1_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableG = SpriteTableG_1_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableG = SpriteTableG_1_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableG = SpriteTableG_1_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_1_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableG = SpriteTableG_1_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableG = SpriteTableG_1_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableG = SpriteTableG_1_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableG = SpriteTableG_1_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableG = SpriteTableG_1_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableG = SpriteTableG_1_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableG = SpriteTableG_1_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableG = SpriteTableG_1_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableG = SpriteTableG_1_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableG = SpriteTableG_1_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableG = SpriteTableG_1_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableG = SpriteTableG_1_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableG = SpriteTableG_1_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableG = SpriteTableG_1_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableG = SpriteTableG_1_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableG = SpriteTableG_1_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableG = SpriteTableG_1_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableG = SpriteTableG_1_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableG = SpriteTableG_1_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableG = SpriteTableG_1_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableG = SpriteTableG_1_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableG = SpriteTableG_1_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableG = SpriteTableG_2_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableG = SpriteTableG_2_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableG = SpriteTableG_2_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableG = SpriteTableG_2_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableG = SpriteTableG_2_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableG = SpriteTableG_2_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableG = SpriteTableG_2_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableG = SpriteTableG_2_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableG = SpriteTableG_2_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableG = SpriteTableG_2_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableG = SpriteTableG_2_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableG = SpriteTableG_2_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableG = SpriteTableG_2_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_2_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableG = SpriteTableG_2_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableG = SpriteTableG_2_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableG = SpriteTableG_2_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableG = SpriteTableG_2_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableG = SpriteTableG_2_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableG = SpriteTableG_2_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableG = SpriteTableG_2_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableG = SpriteTableG_2_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableG = SpriteTableG_2_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableG = SpriteTableG_2_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableG = SpriteTableG_2_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableG = SpriteTableG_2_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableG = SpriteTableG_2_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableG = SpriteTableG_2_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableG = SpriteTableG_2_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableG = SpriteTableG_2_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableG = SpriteTableG_2_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableG = SpriteTableG_2_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableG = SpriteTableG_2_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableG = SpriteTableG_2_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableG = SpriteTableG_2_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableG = SpriteTableG_2_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableG = SpriteTableG_3_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableG = SpriteTableG_3_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableG = SpriteTableG_3_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableG = SpriteTableG_3_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableG = SpriteTableG_3_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableG = SpriteTableG_3_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableG = SpriteTableG_3_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableG = SpriteTableG_3_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableG = SpriteTableG_3_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableG = SpriteTableG_3_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableG = SpriteTableG_3_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableG = SpriteTableG_3_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableG = SpriteTableG_3_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_3_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableG = SpriteTableG_3_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableG = SpriteTableG_3_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableG = SpriteTableG_3_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableG = SpriteTableG_3_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableG = SpriteTableG_3_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableG = SpriteTableG_3_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableG = SpriteTableG_3_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableG = SpriteTableG_3_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableG = SpriteTableG_3_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableG = SpriteTableG_3_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableG = SpriteTableG_3_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableG = SpriteTableG_3_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableG = SpriteTableG_3_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableG = SpriteTableG_3_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableG = SpriteTableG_3_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableG = SpriteTableG_3_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableG = SpriteTableG_3_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableG = SpriteTableG_3_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableG = SpriteTableG_3_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableG = SpriteTableG_3_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableG = SpriteTableG_3_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableG = SpriteTableG_3_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableG = SpriteTableG_4_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableG = SpriteTableG_4_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableG = SpriteTableG_4_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableG = SpriteTableG_4_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableG = SpriteTableG_4_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableG = SpriteTableG_4_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableG = SpriteTableG_4_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableG = SpriteTableG_4_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableG = SpriteTableG_4_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableG = SpriteTableG_4_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableG = SpriteTableG_4_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableG = SpriteTableG_4_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableG = SpriteTableG_4_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_4_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableG = SpriteTableG_4_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableG = SpriteTableG_4_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableG = SpriteTableG_4_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableG = SpriteTableG_4_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableG = SpriteTableG_4_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableG = SpriteTableG_4_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableG = SpriteTableG_4_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableG = SpriteTableG_4_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableG = SpriteTableG_4_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableG = SpriteTableG_4_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableG = SpriteTableG_4_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableG = SpriteTableG_4_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableG = SpriteTableG_4_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableG = SpriteTableG_4_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableG = SpriteTableG_4_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableG = SpriteTableG_4_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableG = SpriteTableG_4_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableG = SpriteTableG_4_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableG = SpriteTableG_4_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableG = SpriteTableG_4_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableG = SpriteTableG_4_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableG = SpriteTableG_4_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableG = SpriteTableG_5_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableG = SpriteTableG_5_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableG = SpriteTableG_5_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableG = SpriteTableG_5_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableG = SpriteTableG_5_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableG = SpriteTableG_5_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableG = SpriteTableG_5_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableG = SpriteTableG_5_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableG = SpriteTableG_5_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableG = SpriteTableG_5_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableG = SpriteTableG_5_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableG = SpriteTableG_5_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableG = SpriteTableG_5_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_5_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableG = SpriteTableG_5_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableG = SpriteTableG_5_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableG = SpriteTableG_5_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableG = SpriteTableG_5_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableG = SpriteTableG_5_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableG = SpriteTableG_5_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableG = SpriteTableG_5_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableG = SpriteTableG_5_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableG = SpriteTableG_5_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableG = SpriteTableG_5_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableG = SpriteTableG_5_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableG = SpriteTableG_5_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableG = SpriteTableG_5_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableG = SpriteTableG_5_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableG = SpriteTableG_5_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableG = SpriteTableG_5_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableG = SpriteTableG_5_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableG = SpriteTableG_5_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableG = SpriteTableG_5_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableG = SpriteTableG_5_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableG = SpriteTableG_5_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableG = SpriteTableG_5_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableG = SpriteTableG_6_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableG = SpriteTableG_6_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableG = SpriteTableG_6_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableG = SpriteTableG_6_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableG = SpriteTableG_6_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableG = SpriteTableG_6_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableG = SpriteTableG_6_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableG = SpriteTableG_6_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableG = SpriteTableG_6_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableG = SpriteTableG_6_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableG = SpriteTableG_6_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableG = SpriteTableG_6_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableG = SpriteTableG_6_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_6_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableG = SpriteTableG_6_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableG = SpriteTableG_6_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableG = SpriteTableG_6_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableG = SpriteTableG_6_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableG = SpriteTableG_6_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableG = SpriteTableG_6_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableG = SpriteTableG_6_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableG = SpriteTableG_6_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableG = SpriteTableG_6_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableG = SpriteTableG_6_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableG = SpriteTableG_6_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableG = SpriteTableG_6_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableG = SpriteTableG_6_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableG = SpriteTableG_6_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableG = SpriteTableG_6_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableG = SpriteTableG_6_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableG = SpriteTableG_6_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableG = SpriteTableG_6_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableG = SpriteTableG_6_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableG = SpriteTableG_6_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableG = SpriteTableG_6_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableG = SpriteTableG_6_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableG = SpriteTableG_7_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableG = SpriteTableG_7_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableG = SpriteTableG_7_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableG = SpriteTableG_7_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableG = SpriteTableG_7_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableG = SpriteTableG_7_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableG = SpriteTableG_7_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableG = SpriteTableG_7_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableG = SpriteTableG_7_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableG = SpriteTableG_7_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableG = SpriteTableG_7_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableG = SpriteTableG_7_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableG = SpriteTableG_7_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_7_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableG = SpriteTableG_7_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableG = SpriteTableG_7_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableG = SpriteTableG_7_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableG = SpriteTableG_7_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableG = SpriteTableG_7_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableG = SpriteTableG_7_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableG = SpriteTableG_7_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableG = SpriteTableG_7_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableG = SpriteTableG_7_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableG = SpriteTableG_7_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableG = SpriteTableG_7_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableG = SpriteTableG_7_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableG = SpriteTableG_7_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableG = SpriteTableG_7_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableG = SpriteTableG_7_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableG = SpriteTableG_7_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableG = SpriteTableG_7_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableG = SpriteTableG_7_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableG = SpriteTableG_7_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableG = SpriteTableG_7_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableG = SpriteTableG_7_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableG = SpriteTableG_7_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableG = SpriteTableG_8_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableG = SpriteTableG_8_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableG = SpriteTableG_8_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableG = SpriteTableG_8_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableG = SpriteTableG_8_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableG = SpriteTableG_8_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableG = SpriteTableG_8_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableG = SpriteTableG_8_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableG = SpriteTableG_8_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableG = SpriteTableG_8_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableG = SpriteTableG_8_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableG = SpriteTableG_8_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableG = SpriteTableG_8_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_8_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableG = SpriteTableG_8_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableG = SpriteTableG_8_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableG = SpriteTableG_8_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableG = SpriteTableG_8_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableG = SpriteTableG_8_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableG = SpriteTableG_8_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableG = SpriteTableG_8_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableG = SpriteTableG_8_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableG = SpriteTableG_8_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableG = SpriteTableG_8_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableG = SpriteTableG_8_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableG = SpriteTableG_8_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableG = SpriteTableG_8_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableG = SpriteTableG_8_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableG = SpriteTableG_8_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableG = SpriteTableG_8_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableG = SpriteTableG_8_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableG = SpriteTableG_8_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableG = SpriteTableG_8_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableG = SpriteTableG_8_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableG = SpriteTableG_8_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableG = SpriteTableG_8_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableG = SpriteTableG_9_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableG = SpriteTableG_9_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableG = SpriteTableG_9_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableG = SpriteTableG_9_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableG = SpriteTableG_9_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableG = SpriteTableG_9_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableG = SpriteTableG_9_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableG = SpriteTableG_9_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableG = SpriteTableG_9_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableG = SpriteTableG_9_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableG = SpriteTableG_9_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableG = SpriteTableG_9_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableG = SpriteTableG_9_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_9_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableG = SpriteTableG_9_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableG = SpriteTableG_9_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableG = SpriteTableG_9_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableG = SpriteTableG_9_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableG = SpriteTableG_9_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableG = SpriteTableG_9_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableG = SpriteTableG_9_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableG = SpriteTableG_9_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableG = SpriteTableG_9_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableG = SpriteTableG_9_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableG = SpriteTableG_9_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableG = SpriteTableG_9_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableG = SpriteTableG_9_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableG = SpriteTableG_9_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableG = SpriteTableG_9_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableG = SpriteTableG_9_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableG = SpriteTableG_9_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableG = SpriteTableG_9_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableG = SpriteTableG_9_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableG = SpriteTableG_9_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableG = SpriteTableG_9_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableG = SpriteTableG_9_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableG = SpriteTableG_10_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableG = SpriteTableG_10_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableG = SpriteTableG_10_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableG = SpriteTableG_10_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableG = SpriteTableG_10_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableG = SpriteTableG_10_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableG = SpriteTableG_10_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableG = SpriteTableG_10_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableG = SpriteTableG_10_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableG = SpriteTableG_10_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableG = SpriteTableG_10_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableG = SpriteTableG_10_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableG = SpriteTableG_10_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_10_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableG = SpriteTableG_10_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableG = SpriteTableG_10_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableG = SpriteTableG_10_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableG = SpriteTableG_10_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableG = SpriteTableG_10_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableG = SpriteTableG_10_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableG = SpriteTableG_10_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableG = SpriteTableG_10_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableG = SpriteTableG_10_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableG = SpriteTableG_10_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableG = SpriteTableG_10_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableG = SpriteTableG_10_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableG = SpriteTableG_10_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableG = SpriteTableG_10_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableG = SpriteTableG_10_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableG = SpriteTableG_10_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableG = SpriteTableG_10_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableG = SpriteTableG_10_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableG = SpriteTableG_10_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableG = SpriteTableG_10_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableG = SpriteTableG_10_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableG = SpriteTableG_10_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableG = SpriteTableG_11_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableG = SpriteTableG_11_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableG = SpriteTableG_11_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableG = SpriteTableG_11_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableG = SpriteTableG_11_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableG = SpriteTableG_11_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableG = SpriteTableG_11_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableG = SpriteTableG_11_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableG = SpriteTableG_11_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableG = SpriteTableG_11_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableG = SpriteTableG_11_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableG = SpriteTableG_11_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableG = SpriteTableG_11_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_11_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableG = SpriteTableG_11_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableG = SpriteTableG_11_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableG = SpriteTableG_11_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableG = SpriteTableG_11_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableG = SpriteTableG_11_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableG = SpriteTableG_11_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableG = SpriteTableG_11_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableG = SpriteTableG_11_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableG = SpriteTableG_11_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableG = SpriteTableG_11_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableG = SpriteTableG_11_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableG = SpriteTableG_11_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableG = SpriteTableG_11_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableG = SpriteTableG_11_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableG = SpriteTableG_11_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableG = SpriteTableG_11_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableG = SpriteTableG_11_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableG = SpriteTableG_11_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableG = SpriteTableG_11_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableG = SpriteTableG_11_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableG = SpriteTableG_11_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableG = SpriteTableG_11_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableG = SpriteTableG_12_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableG = SpriteTableG_12_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableG = SpriteTableG_12_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableG = SpriteTableG_12_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableG = SpriteTableG_12_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableG = SpriteTableG_12_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableG = SpriteTableG_12_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableG = SpriteTableG_12_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableG = SpriteTableG_12_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableG = SpriteTableG_12_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableG = SpriteTableG_12_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableG = SpriteTableG_12_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableG = SpriteTableG_12_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_12_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableG = SpriteTableG_12_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableG = SpriteTableG_12_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableG = SpriteTableG_12_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableG = SpriteTableG_12_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableG = SpriteTableG_12_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableG = SpriteTableG_12_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableG = SpriteTableG_12_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableG = SpriteTableG_12_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableG = SpriteTableG_12_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableG = SpriteTableG_12_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableG = SpriteTableG_12_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableG = SpriteTableG_12_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableG = SpriteTableG_12_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableG = SpriteTableG_12_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableG = SpriteTableG_12_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableG = SpriteTableG_12_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableG = SpriteTableG_12_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableG = SpriteTableG_12_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableG = SpriteTableG_12_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableG = SpriteTableG_12_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableG = SpriteTableG_12_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableG = SpriteTableG_12_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableG = SpriteTableG_13_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableG = SpriteTableG_13_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableG = SpriteTableG_13_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableG = SpriteTableG_13_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableG = SpriteTableG_13_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableG = SpriteTableG_13_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableG = SpriteTableG_13_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableG = SpriteTableG_13_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableG = SpriteTableG_13_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableG = SpriteTableG_13_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableG = SpriteTableG_13_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableG = SpriteTableG_13_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableG = SpriteTableG_13_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_13_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableG = SpriteTableG_13_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableG = SpriteTableG_13_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableG = SpriteTableG_13_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableG = SpriteTableG_13_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableG = SpriteTableG_13_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableG = SpriteTableG_13_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableG = SpriteTableG_13_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableG = SpriteTableG_13_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableG = SpriteTableG_13_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableG = SpriteTableG_13_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableG = SpriteTableG_13_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableG = SpriteTableG_13_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableG = SpriteTableG_13_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableG = SpriteTableG_13_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableG = SpriteTableG_13_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableG = SpriteTableG_13_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableG = SpriteTableG_13_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableG = SpriteTableG_13_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableG = SpriteTableG_13_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableG = SpriteTableG_13_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableG = SpriteTableG_13_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableG = SpriteTableG_13_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableG = SpriteTableG_14_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableG = SpriteTableG_14_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableG = SpriteTableG_14_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableG = SpriteTableG_14_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableG = SpriteTableG_14_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableG = SpriteTableG_14_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableG = SpriteTableG_14_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableG = SpriteTableG_14_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableG = SpriteTableG_14_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableG = SpriteTableG_14_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableG = SpriteTableG_14_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableG = SpriteTableG_14_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableG = SpriteTableG_14_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_14_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableG = SpriteTableG_14_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableG = SpriteTableG_14_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableG = SpriteTableG_14_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableG = SpriteTableG_14_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableG = SpriteTableG_14_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableG = SpriteTableG_14_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableG = SpriteTableG_14_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableG = SpriteTableG_14_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableG = SpriteTableG_14_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableG = SpriteTableG_14_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableG = SpriteTableG_14_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableG = SpriteTableG_14_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableG = SpriteTableG_14_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableG = SpriteTableG_14_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableG = SpriteTableG_14_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableG = SpriteTableG_14_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableG = SpriteTableG_14_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableG = SpriteTableG_14_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableG = SpriteTableG_14_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableG = SpriteTableG_14_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableG = SpriteTableG_14_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableG = SpriteTableG_14_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableG = SpriteTableG_15_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableG = SpriteTableG_15_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableG = SpriteTableG_15_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableG = SpriteTableG_15_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableG = SpriteTableG_15_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableG = SpriteTableG_15_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableG = SpriteTableG_15_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableG = SpriteTableG_15_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableG = SpriteTableG_15_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableG = SpriteTableG_15_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableG = SpriteTableG_15_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableG = SpriteTableG_15_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableG = SpriteTableG_15_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_15_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableG = SpriteTableG_15_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableG = SpriteTableG_15_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableG = SpriteTableG_15_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableG = SpriteTableG_15_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableG = SpriteTableG_15_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableG = SpriteTableG_15_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableG = SpriteTableG_15_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableG = SpriteTableG_15_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableG = SpriteTableG_15_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableG = SpriteTableG_15_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableG = SpriteTableG_15_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableG = SpriteTableG_15_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableG = SpriteTableG_15_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableG = SpriteTableG_15_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableG = SpriteTableG_15_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableG = SpriteTableG_15_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableG = SpriteTableG_15_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableG = SpriteTableG_15_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableG = SpriteTableG_15_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableG = SpriteTableG_15_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableG = SpriteTableG_15_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableG = SpriteTableG_15_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableG = SpriteTableG_16_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableG = SpriteTableG_16_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableG = SpriteTableG_16_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableG = SpriteTableG_16_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableG = SpriteTableG_16_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableG = SpriteTableG_16_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableG = SpriteTableG_16_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableG = SpriteTableG_16_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableG = SpriteTableG_16_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableG = SpriteTableG_16_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableG = SpriteTableG_16_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableG = SpriteTableG_16_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableG = SpriteTableG_16_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_16_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableG = SpriteTableG_16_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableG = SpriteTableG_16_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableG = SpriteTableG_16_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableG = SpriteTableG_16_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableG = SpriteTableG_16_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableG = SpriteTableG_16_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableG = SpriteTableG_16_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableG = SpriteTableG_16_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableG = SpriteTableG_16_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableG = SpriteTableG_16_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableG = SpriteTableG_16_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableG = SpriteTableG_16_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableG = SpriteTableG_16_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableG = SpriteTableG_16_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableG = SpriteTableG_16_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableG = SpriteTableG_16_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableG = SpriteTableG_16_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableG = SpriteTableG_16_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableG = SpriteTableG_16_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableG = SpriteTableG_16_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableG = SpriteTableG_16_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableG = SpriteTableG_16_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableG = SpriteTableG_17_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableG = SpriteTableG_17_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableG = SpriteTableG_17_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableG = SpriteTableG_17_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableG = SpriteTableG_17_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableG = SpriteTableG_17_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableG = SpriteTableG_17_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableG = SpriteTableG_17_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableG = SpriteTableG_17_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableG = SpriteTableG_17_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableG = SpriteTableG_17_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableG = SpriteTableG_17_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableG = SpriteTableG_17_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_17_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableG = SpriteTableG_17_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableG = SpriteTableG_17_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableG = SpriteTableG_17_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableG = SpriteTableG_17_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableG = SpriteTableG_17_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableG = SpriteTableG_17_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableG = SpriteTableG_17_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableG = SpriteTableG_17_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableG = SpriteTableG_17_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableG = SpriteTableG_17_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableG = SpriteTableG_17_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableG = SpriteTableG_17_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableG = SpriteTableG_17_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableG = SpriteTableG_17_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableG = SpriteTableG_17_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableG = SpriteTableG_17_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableG = SpriteTableG_17_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableG = SpriteTableG_17_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableG = SpriteTableG_17_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableG = SpriteTableG_17_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableG = SpriteTableG_17_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableG = SpriteTableG_17_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableG = SpriteTableG_18_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableG = SpriteTableG_18_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableG = SpriteTableG_18_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableG = SpriteTableG_18_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableG = SpriteTableG_18_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableG = SpriteTableG_18_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableG = SpriteTableG_18_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableG = SpriteTableG_18_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableG = SpriteTableG_18_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableG = SpriteTableG_18_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableG = SpriteTableG_18_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableG = SpriteTableG_18_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableG = SpriteTableG_18_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_18_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableG = SpriteTableG_18_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableG = SpriteTableG_18_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableG = SpriteTableG_18_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableG = SpriteTableG_18_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableG = SpriteTableG_18_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableG = SpriteTableG_18_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableG = SpriteTableG_18_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableG = SpriteTableG_18_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableG = SpriteTableG_18_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableG = SpriteTableG_18_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableG = SpriteTableG_18_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableG = SpriteTableG_18_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableG = SpriteTableG_18_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableG = SpriteTableG_18_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableG = SpriteTableG_18_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableG = SpriteTableG_18_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableG = SpriteTableG_18_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableG = SpriteTableG_18_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableG = SpriteTableG_18_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableG = SpriteTableG_18_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableG = SpriteTableG_18_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableG = SpriteTableG_18_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableG = SpriteTableG_19_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableG = SpriteTableG_19_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableG = SpriteTableG_19_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableG = SpriteTableG_19_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableG = SpriteTableG_19_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableG = SpriteTableG_19_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableG = SpriteTableG_19_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableG = SpriteTableG_19_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableG = SpriteTableG_19_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableG = SpriteTableG_19_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableG = SpriteTableG_19_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableG = SpriteTableG_19_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableG = SpriteTableG_19_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_19_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableG = SpriteTableG_19_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableG = SpriteTableG_19_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableG = SpriteTableG_19_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableG = SpriteTableG_19_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableG = SpriteTableG_19_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableG = SpriteTableG_19_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableG = SpriteTableG_19_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableG = SpriteTableG_19_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableG = SpriteTableG_19_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableG = SpriteTableG_19_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableG = SpriteTableG_19_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableG = SpriteTableG_19_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableG = SpriteTableG_19_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableG = SpriteTableG_19_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableG = SpriteTableG_19_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableG = SpriteTableG_19_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableG = SpriteTableG_19_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableG = SpriteTableG_19_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableG = SpriteTableG_19_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableG = SpriteTableG_19_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableG = SpriteTableG_19_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableG = SpriteTableG_19_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableG = SpriteTableG_20_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableG = SpriteTableG_20_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableG = SpriteTableG_20_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableG = SpriteTableG_20_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableG = SpriteTableG_20_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableG = SpriteTableG_20_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableG = SpriteTableG_20_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableG = SpriteTableG_20_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableG = SpriteTableG_20_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableG = SpriteTableG_20_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableG = SpriteTableG_20_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableG = SpriteTableG_20_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableG = SpriteTableG_20_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_20_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableG = SpriteTableG_20_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableG = SpriteTableG_20_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableG = SpriteTableG_20_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableG = SpriteTableG_20_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableG = SpriteTableG_20_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableG = SpriteTableG_20_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableG = SpriteTableG_20_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableG = SpriteTableG_20_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableG = SpriteTableG_20_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableG = SpriteTableG_20_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableG = SpriteTableG_20_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableG = SpriteTableG_20_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableG = SpriteTableG_20_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableG = SpriteTableG_20_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableG = SpriteTableG_20_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableG = SpriteTableG_20_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableG = SpriteTableG_20_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableG = SpriteTableG_20_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableG = SpriteTableG_20_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableG = SpriteTableG_20_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableG = SpriteTableG_20_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableG = SpriteTableG_20_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableG = SpriteTableG_21_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableG = SpriteTableG_21_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableG = SpriteTableG_21_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableG = SpriteTableG_21_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableG = SpriteTableG_21_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableG = SpriteTableG_21_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableG = SpriteTableG_21_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableG = SpriteTableG_21_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableG = SpriteTableG_21_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableG = SpriteTableG_21_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableG = SpriteTableG_21_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableG = SpriteTableG_21_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableG = SpriteTableG_21_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_21_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableG = SpriteTableG_21_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableG = SpriteTableG_21_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableG = SpriteTableG_21_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableG = SpriteTableG_21_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableG = SpriteTableG_21_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableG = SpriteTableG_21_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableG = SpriteTableG_21_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableG = SpriteTableG_21_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableG = SpriteTableG_21_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableG = SpriteTableG_21_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableG = SpriteTableG_21_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableG = SpriteTableG_21_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableG = SpriteTableG_21_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableG = SpriteTableG_21_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableG = SpriteTableG_21_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableG = SpriteTableG_21_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableG = SpriteTableG_21_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableG = SpriteTableG_21_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableG = SpriteTableG_21_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableG = SpriteTableG_21_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableG = SpriteTableG_21_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableG = SpriteTableG_21_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableG = SpriteTableG_22_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableG = SpriteTableG_22_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableG = SpriteTableG_22_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableG = SpriteTableG_22_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableG = SpriteTableG_22_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableG = SpriteTableG_22_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableG = SpriteTableG_22_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableG = SpriteTableG_22_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableG = SpriteTableG_22_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableG = SpriteTableG_22_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableG = SpriteTableG_22_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableG = SpriteTableG_22_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableG = SpriteTableG_22_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_22_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableG = SpriteTableG_22_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableG = SpriteTableG_22_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableG = SpriteTableG_22_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableG = SpriteTableG_22_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableG = SpriteTableG_22_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableG = SpriteTableG_22_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableG = SpriteTableG_22_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableG = SpriteTableG_22_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableG = SpriteTableG_22_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableG = SpriteTableG_22_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableG = SpriteTableG_22_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableG = SpriteTableG_22_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableG = SpriteTableG_22_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableG = SpriteTableG_22_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableG = SpriteTableG_22_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableG = SpriteTableG_22_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableG = SpriteTableG_22_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableG = SpriteTableG_22_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableG = SpriteTableG_22_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableG = SpriteTableG_22_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableG = SpriteTableG_22_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableG = SpriteTableG_22_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableG = SpriteTableG_23_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableG = SpriteTableG_23_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableG = SpriteTableG_23_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableG = SpriteTableG_23_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableG = SpriteTableG_23_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableG = SpriteTableG_23_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableG = SpriteTableG_23_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableG = SpriteTableG_23_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableG = SpriteTableG_23_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableG = SpriteTableG_23_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableG = SpriteTableG_23_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableG = SpriteTableG_23_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableG = SpriteTableG_23_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_23_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableG = SpriteTableG_23_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableG = SpriteTableG_23_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableG = SpriteTableG_23_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableG = SpriteTableG_23_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableG = SpriteTableG_23_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableG = SpriteTableG_23_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableG = SpriteTableG_23_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableG = SpriteTableG_23_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableG = SpriteTableG_23_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableG = SpriteTableG_23_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableG = SpriteTableG_23_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableG = SpriteTableG_23_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableG = SpriteTableG_23_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableG = SpriteTableG_23_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableG = SpriteTableG_23_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableG = SpriteTableG_23_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableG = SpriteTableG_23_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableG = SpriteTableG_23_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableG = SpriteTableG_23_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableG = SpriteTableG_23_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableG = SpriteTableG_23_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableG = SpriteTableG_23_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableG = SpriteTableG_24_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableG = SpriteTableG_24_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableG = SpriteTableG_24_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableG = SpriteTableG_24_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableG = SpriteTableG_24_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableG = SpriteTableG_24_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableG = SpriteTableG_24_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableG = SpriteTableG_24_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableG = SpriteTableG_24_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableG = SpriteTableG_24_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableG = SpriteTableG_24_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableG = SpriteTableG_24_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableG = SpriteTableG_24_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_24_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableG = SpriteTableG_24_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableG = SpriteTableG_24_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableG = SpriteTableG_24_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableG = SpriteTableG_24_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableG = SpriteTableG_24_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableG = SpriteTableG_24_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableG = SpriteTableG_24_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableG = SpriteTableG_24_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableG = SpriteTableG_24_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableG = SpriteTableG_24_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableG = SpriteTableG_24_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableG = SpriteTableG_24_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableG = SpriteTableG_24_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableG = SpriteTableG_24_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableG = SpriteTableG_24_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableG = SpriteTableG_24_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableG = SpriteTableG_24_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableG = SpriteTableG_24_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableG = SpriteTableG_24_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableG = SpriteTableG_24_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableG = SpriteTableG_24_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableG = SpriteTableG_24_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableG = SpriteTableG_25_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableG = SpriteTableG_25_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableG = SpriteTableG_25_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableG = SpriteTableG_25_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableG = SpriteTableG_25_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableG = SpriteTableG_25_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableG = SpriteTableG_25_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableG = SpriteTableG_25_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableG = SpriteTableG_25_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableG = SpriteTableG_25_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableG = SpriteTableG_25_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableG = SpriteTableG_25_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableG = SpriteTableG_25_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_25_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableG = SpriteTableG_25_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableG = SpriteTableG_25_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableG = SpriteTableG_25_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableG = SpriteTableG_25_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableG = SpriteTableG_25_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableG = SpriteTableG_25_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableG = SpriteTableG_25_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableG = SpriteTableG_25_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableG = SpriteTableG_25_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableG = SpriteTableG_25_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableG = SpriteTableG_25_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableG = SpriteTableG_25_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableG = SpriteTableG_25_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableG = SpriteTableG_25_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableG = SpriteTableG_25_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableG = SpriteTableG_25_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableG = SpriteTableG_25_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableG = SpriteTableG_25_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableG = SpriteTableG_25_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableG = SpriteTableG_25_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableG = SpriteTableG_25_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableG = SpriteTableG_25_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableG = SpriteTableG_26_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableG = SpriteTableG_26_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableG = SpriteTableG_26_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableG = SpriteTableG_26_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableG = SpriteTableG_26_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableG = SpriteTableG_26_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableG = SpriteTableG_26_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableG = SpriteTableG_26_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableG = SpriteTableG_26_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableG = SpriteTableG_26_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableG = SpriteTableG_26_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableG = SpriteTableG_26_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableG = SpriteTableG_26_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_26_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableG = SpriteTableG_26_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableG = SpriteTableG_26_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableG = SpriteTableG_26_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableG = SpriteTableG_26_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableG = SpriteTableG_26_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableG = SpriteTableG_26_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableG = SpriteTableG_26_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableG = SpriteTableG_26_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableG = SpriteTableG_26_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableG = SpriteTableG_26_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableG = SpriteTableG_26_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableG = SpriteTableG_26_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableG = SpriteTableG_26_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableG = SpriteTableG_26_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableG = SpriteTableG_26_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableG = SpriteTableG_26_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableG = SpriteTableG_26_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableG = SpriteTableG_26_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableG = SpriteTableG_26_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableG = SpriteTableG_26_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableG = SpriteTableG_26_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableG = SpriteTableG_26_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableG = SpriteTableG_27_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableG = SpriteTableG_27_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableG = SpriteTableG_27_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableG = SpriteTableG_27_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableG = SpriteTableG_27_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableG = SpriteTableG_27_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableG = SpriteTableG_27_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableG = SpriteTableG_27_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableG = SpriteTableG_27_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableG = SpriteTableG_27_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableG = SpriteTableG_27_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableG = SpriteTableG_27_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableG = SpriteTableG_27_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_27_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableG = SpriteTableG_27_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableG = SpriteTableG_27_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableG = SpriteTableG_27_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableG = SpriteTableG_27_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableG = SpriteTableG_27_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableG = SpriteTableG_27_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableG = SpriteTableG_27_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableG = SpriteTableG_27_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableG = SpriteTableG_27_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableG = SpriteTableG_27_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableG = SpriteTableG_27_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableG = SpriteTableG_27_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableG = SpriteTableG_27_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableG = SpriteTableG_27_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableG = SpriteTableG_27_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableG = SpriteTableG_27_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableG = SpriteTableG_27_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableG = SpriteTableG_27_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableG = SpriteTableG_27_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableG = SpriteTableG_27_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableG = SpriteTableG_27_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableG = SpriteTableG_27_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableG = SpriteTableG_28_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableG = SpriteTableG_28_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableG = SpriteTableG_28_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableG = SpriteTableG_28_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableG = SpriteTableG_28_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableG = SpriteTableG_28_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableG = SpriteTableG_28_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableG = SpriteTableG_28_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableG = SpriteTableG_28_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableG = SpriteTableG_28_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableG = SpriteTableG_28_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableG = SpriteTableG_28_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableG = SpriteTableG_28_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_28_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableG = SpriteTableG_28_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableG = SpriteTableG_28_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableG = SpriteTableG_28_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableG = SpriteTableG_28_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableG = SpriteTableG_28_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableG = SpriteTableG_28_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableG = SpriteTableG_28_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableG = SpriteTableG_28_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableG = SpriteTableG_28_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableG = SpriteTableG_28_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableG = SpriteTableG_28_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableG = SpriteTableG_28_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableG = SpriteTableG_28_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableG = SpriteTableG_28_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableG = SpriteTableG_28_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableG = SpriteTableG_28_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableG = SpriteTableG_28_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableG = SpriteTableG_28_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableG = SpriteTableG_28_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableG = SpriteTableG_28_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableG = SpriteTableG_28_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableG = SpriteTableG_28_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableG = SpriteTableG_29_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableG = SpriteTableG_29_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableG = SpriteTableG_29_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableG = SpriteTableG_29_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableG = SpriteTableG_29_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableG = SpriteTableG_29_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableG = SpriteTableG_29_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableG = SpriteTableG_29_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableG = SpriteTableG_29_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableG = SpriteTableG_29_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableG = SpriteTableG_29_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableG = SpriteTableG_29_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableG = SpriteTableG_29_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_29_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableG = SpriteTableG_29_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableG = SpriteTableG_29_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableG = SpriteTableG_29_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableG = SpriteTableG_29_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableG = SpriteTableG_29_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableG = SpriteTableG_29_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableG = SpriteTableG_29_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableG = SpriteTableG_29_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableG = SpriteTableG_29_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableG = SpriteTableG_29_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableG = SpriteTableG_29_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableG = SpriteTableG_29_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableG = SpriteTableG_29_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableG = SpriteTableG_29_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableG = SpriteTableG_29_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableG = SpriteTableG_29_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableG = SpriteTableG_29_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableG = SpriteTableG_29_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableG = SpriteTableG_29_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableG = SpriteTableG_29_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableG = SpriteTableG_29_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableG = SpriteTableG_29_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableG = SpriteTableG_30_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableG = SpriteTableG_30_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableG = SpriteTableG_30_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableG = SpriteTableG_30_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableG = SpriteTableG_30_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableG = SpriteTableG_30_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableG = SpriteTableG_30_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableG = SpriteTableG_30_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableG = SpriteTableG_30_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableG = SpriteTableG_30_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableG = SpriteTableG_30_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableG = SpriteTableG_30_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableG = SpriteTableG_30_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_30_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableG = SpriteTableG_30_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableG = SpriteTableG_30_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableG = SpriteTableG_30_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableG = SpriteTableG_30_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableG = SpriteTableG_30_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableG = SpriteTableG_30_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableG = SpriteTableG_30_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableG = SpriteTableG_30_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableG = SpriteTableG_30_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableG = SpriteTableG_30_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableG = SpriteTableG_30_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableG = SpriteTableG_30_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableG = SpriteTableG_30_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableG = SpriteTableG_30_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableG = SpriteTableG_30_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableG = SpriteTableG_30_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableG = SpriteTableG_30_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableG = SpriteTableG_30_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableG = SpriteTableG_30_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableG = SpriteTableG_30_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableG = SpriteTableG_30_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableG = SpriteTableG_30_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableG = SpriteTableG_31_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableG = SpriteTableG_31_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableG = SpriteTableG_31_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableG = SpriteTableG_31_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableG = SpriteTableG_31_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableG = SpriteTableG_31_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableG = SpriteTableG_31_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableG = SpriteTableG_31_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableG = SpriteTableG_31_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableG = SpriteTableG_31_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableG = SpriteTableG_31_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableG = SpriteTableG_31_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableG = SpriteTableG_31_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableG = SpriteTableG_31_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableG = SpriteTableG_31_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableG = SpriteTableG_31_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableG = SpriteTableG_31_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableG = SpriteTableG_31_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableG = SpriteTableG_31_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableG = SpriteTableG_31_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableG = SpriteTableG_31_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableG = SpriteTableG_31_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableG = SpriteTableG_31_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableG = SpriteTableG_31_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableG = SpriteTableG_31_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableG = SpriteTableG_31_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableG = SpriteTableG_31_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableG = SpriteTableG_31_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableG = SpriteTableG_31_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableG = SpriteTableG_31_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableG = SpriteTableG_31_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableG = SpriteTableG_31_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableG = SpriteTableG_31_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableG = SpriteTableG_31_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableG = SpriteTableG_31_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableG = SpriteTableG_31_35[Y_Index][X_Index];
		end
	end

parameter bit [2:0] SpriteTableG_0_0[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_0_1[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_0_2[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_0_3[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_0_4[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_0_5[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_0_6[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd1}};

parameter bit [2:0] SpriteTableG_0_7[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd3,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0}};

parameter bit [2:0] SpriteTableG_0_8[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd4,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd3,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2}};

parameter bit [2:0] SpriteTableG_0_9[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd1}};

parameter bit [2:0] SpriteTableG_0_10[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2,3'd1},
'{3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd1},
'{3'd0,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1},
'{3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1},
'{3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_0_11[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_0_12[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_0_13[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_0_14[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_0_15[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_0_16[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_0_17[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_0_18[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0}};

parameter bit [2:0] SpriteTableG_0_19[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_0_20[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_0_21[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_0_22[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_0_23[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1}};

parameter bit [2:0] SpriteTableG_0_24[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_0_25[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_0_26[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd1},
'{3'd0,3'd0,3'd0,3'd1,3'd2,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd2,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3}};

parameter bit [2:0] SpriteTableG_0_27[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_0_28[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_0_29[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_0_30[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_0_31[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_0_32[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_0_33[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_0_34[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableG_0_35[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_1_0[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_1_1[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_1_2[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_1_3[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_1_4[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd4,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_1_5[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd4,3'd3,3'd1,3'd1,3'd3,3'd4,3'd1},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd4,3'd1},
'{3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd4,3'd4,3'd4,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_1_6[7:0][7:0] = '{'{3'd0,3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_1_7[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd4,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_1_8[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd1,3'd0,3'd0},
'{3'd1,3'd4,3'd4,3'd1,3'd1,3'd4,3'd0,3'd0},
'{3'd2,3'd2,3'd2,3'd3,3'd1,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_1_9[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd2,3'd1,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd3,3'd4,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd3,3'd1,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd2,3'd3,3'd1,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd3,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd3},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1}};

parameter bit [2:0] SpriteTableG_1_10[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1}};

parameter bit [2:0] SpriteTableG_1_11[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_1_12[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_1_13[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_1_14[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_1_15[7:0][7:0] = '{'{3'd0,3'd4,3'd2,3'd3,3'd2,3'd0,3'd1,3'd0},
'{3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd2,3'd3,3'd3,3'd3,3'd2},
'{3'd0,3'd0,3'd0,3'd4,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd4,3'd3,3'd2,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd4,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_1_16[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_1_17[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd3,3'd2,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd2,3'd3,3'd2,3'd0,3'd0,3'd0},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd1},
'{3'd1,3'd2,3'd2,3'd3,3'd3,3'd2,3'd2,3'd2},
'{3'd0,3'd2,3'd2,3'd3,3'd3,3'd2,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_1_18[7:0][7:0] = '{'{3'd0,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0},
'{3'd4,3'd3,3'd2,3'd1,3'd3,3'd2,3'd0,3'd0},
'{3'd4,3'd1,3'd0,3'd0,3'd1,3'd1,3'd0,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0},
'{3'd0,3'd0,3'd1,3'd1,3'd0,3'd1,3'd1,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_1_19[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd2},
'{3'd1,3'd1,3'd4,3'd0,3'd1,3'd1,3'd0,3'd1},
'{3'd2,3'd2,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0}};

parameter bit [2:0] SpriteTableG_1_20[7:0][7:0] = '{'{3'd0,3'd1,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd0,3'd1,3'd1,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd1,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1}};

parameter bit [2:0] SpriteTableG_1_21[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_1_22[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1}};

parameter bit [2:0] SpriteTableG_1_23[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd0,3'd1,3'd0,3'd0,3'd0,3'd1},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd2,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_1_24[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0},
'{3'd1,3'd0,3'd1,3'd2,3'd3,3'd3,3'd0,3'd0},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd0},
'{3'd3,3'd3,3'd3,3'd2,3'd2,3'd3,3'd3,3'd1},
'{3'd2,3'd3,3'd2,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd2,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_1_25[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd3}};

parameter bit [2:0] SpriteTableG_1_26[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd4,3'd1,3'd2,3'd3,3'd3},
'{3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_1_27[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_1_28[7:0][7:0] = '{'{3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0},
'{3'd0,3'd2,3'd3,3'd2,3'd4,3'd0,3'd0,3'd0},
'{3'd0,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_1_29[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_1_30[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3}};

parameter bit [2:0] SpriteTableG_1_31[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd3,3'd4},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd0,3'd0,3'd0,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd0,3'd0,3'd0,3'd1,3'd3,3'd2,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd1,3'd3,3'd2,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_1_32[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd2,3'd3,3'd2,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd1,3'd2,3'd4,3'd1,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_1_33[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd0,3'd0,3'd0,3'd4,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_1_34[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableG_1_35[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_2_0[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_2_1[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_2_2[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_2_3[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_2_4[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd4,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_2_5[7:0][7:0] = '{'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd1,3'd1,3'd1},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd3,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3}};

parameter bit [2:0] SpriteTableG_2_6[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1}};

parameter bit [2:0] SpriteTableG_2_7[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd0,3'd0,3'd4,3'd1,3'd4,3'd4,3'd1,3'd3},
'{3'd0,3'd0,3'd0,3'd4,3'd1,3'd1,3'd1,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_2_8[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_2_9[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd2},
'{3'd3,3'd1,3'd1,3'd1,3'd3,3'd3,3'd2,3'd1},
'{3'd2,3'd2,3'd3,3'd2,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1}};

parameter bit [2:0] SpriteTableG_2_10[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_2_11[7:0][7:0] = '{'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_2_12[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd4,3'd4,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd3,3'd1,3'd4,3'd2,3'd2},
'{3'd0,3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd0,3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd4},
'{3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd0,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_2_13[7:0][7:0] = '{'{3'd0,3'd4,3'd4,3'd2,3'd3,3'd3,3'd2,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd3,3'd2,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd2,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_2_14[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_2_15[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd0,3'd1,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd1,3'd0,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd2,3'd0,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd1}};

parameter bit [2:0] SpriteTableG_2_16[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd4,3'd3,3'd4,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd4,3'd1,3'd4,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_2_17[7:0][7:0] = '{'{3'd1,3'd0,3'd0,3'd4,3'd3,3'd4,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd4,3'd3,3'd4,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd4,3'd0,3'd0,3'd4,3'd3,3'd4,3'd0,3'd1},
'{3'd1,3'd0,3'd0,3'd1,3'd3,3'd2,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_2_18[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd1,3'd0},
'{3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2},
'{3'd1,3'd0,3'd0,3'd1,3'd2,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_2_19[7:0][7:0] = '{'{3'd1,3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd1,3'd0,3'd1,3'd2,3'd2,3'd3,3'd3},
'{3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0},
'{3'd1,3'd0,3'd1,3'd1,3'd0,3'd0,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd1}};

parameter bit [2:0] SpriteTableG_2_20[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd1},
'{3'd1,3'd0,3'd0,3'd1,3'd3,3'd1,3'd0,3'd1},
'{3'd1,3'd0,3'd0,3'd1,3'd3,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd1,3'd1,3'd1},
'{3'd1,3'd0,3'd0,3'd1,3'd3,3'd2,3'd1,3'd2}};

parameter bit [2:0] SpriteTableG_2_21[7:0][7:0] = '{'{3'd1,3'd0,3'd0,3'd1,3'd3,3'd2,3'd2,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd4,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd4,3'd3,3'd4,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd1,3'd3,3'd1,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0}};

parameter bit [2:0] SpriteTableG_2_22[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd1},
'{3'd4,3'd0,3'd0,3'd4,3'd2,3'd0,3'd0,3'd1},
'{3'd1,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd1}};

parameter bit [2:0] SpriteTableG_2_23[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd3},
'{3'd0,3'd0,3'd0,3'd1,3'd0,3'd2,3'd3,3'd3},
'{3'd1,3'd0,3'd1,3'd0,3'd2,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd0,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd2,3'd1,3'd1},
'{3'd0,3'd2,3'd2,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_2_24[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_2_25[7:0][7:0] = '{'{3'd0,3'd3,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd3,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_2_26[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_2_27[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_2_28[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd0,3'd0,3'd4,3'd2,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd1,3'd1,3'd1,3'd4,3'd1,3'd3,3'd3,3'd2},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_2_29[7:0][7:0] = '{'{3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd2,3'd2,3'd1,3'd0,3'd2,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd1},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd4,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_2_30[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd4,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd4,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd3,3'd1,3'd1,3'd4,3'd0,3'd4,3'd0},
'{3'd3,3'd1,3'd0,3'd0,3'd4,3'd1,3'd1,3'd1},
'{3'd1,3'd0,3'd0,3'd0,3'd4,3'd4,3'd0,3'd4}};

parameter bit [2:0] SpriteTableG_2_31[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd0},
'{3'd3,3'd4,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0}};

parameter bit [2:0] SpriteTableG_2_32[7:0][7:0] = '{'{3'd3,3'd1,3'd1,3'd4,3'd4,3'd1,3'd1,3'd0},
'{3'd2,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd4},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_2_33[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2}};

parameter bit [2:0] SpriteTableG_2_34[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd4,3'd4,3'd4,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_2_35[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd4,3'd0,3'd0,3'd0},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd0,3'd0,3'd0},
'{3'd4,3'd4,3'd4,3'd1,3'd4,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd4,3'd0,3'd0,3'd0},
'{3'd4,3'd4,3'd4,3'd4,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_3_0[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_3_1[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd3,3'd3,3'd2,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd2,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd2,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_3_2[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd4,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd4,3'd1,3'd4,3'd2,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_3_3[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd3,3'd3,3'd2}};

parameter bit [2:0] SpriteTableG_3_4[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd1,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd4,3'd4},
'{3'd0,3'd0,3'd4,3'd3,3'd1,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_3_5[7:0][7:0] = '{'{3'd1,3'd1,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd0,3'd0,3'd4,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_3_6[7:0][7:0] = '{'{3'd1,3'd0,3'd0,3'd1,3'd4,3'd0,3'd0,3'd0},
'{3'd3,3'd4,3'd0,3'd4,3'd1,3'd0,3'd4,3'd1},
'{3'd1,3'd1,3'd0,3'd0,3'd1,3'd4,3'd4,3'd1},
'{3'd1,3'd1,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0},
'{3'd1,3'd3,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0},
'{3'd1,3'd3,3'd4,3'd0,3'd4,3'd1,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd0,3'd0,3'd3,3'd4,3'd0},
'{3'd4,3'd1,3'd1,3'd0,3'd0,3'd3,3'd4,3'd0}};

parameter bit [2:0] SpriteTableG_3_7[7:0][7:0] = '{'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd3,3'd1,3'd1},
'{3'd0,3'd3,3'd1,3'd0,3'd0,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd0,3'd0,3'd0,3'd3,3'd1,3'd0},
'{3'd3,3'd1,3'd0,3'd0,3'd0,3'd3,3'd4,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd4,3'd3,3'd2,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_3_8[7:0][7:0] = '{'{3'd0,3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2},
'{3'd1,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd1},
'{3'd1,3'd3,3'd2,3'd4,3'd4,3'd1,3'd1,3'd1},
'{3'd1,3'd3,3'd4,3'd0,3'd0,3'd2,3'd1,3'd2},
'{3'd2,3'd2,3'd0,3'd0,3'd4,3'd1,3'd0,3'd1}};

parameter bit [2:0] SpriteTableG_3_9[7:0][7:0] = '{'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_3_10[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_3_11[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_3_12[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0},
'{3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_3_13[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd2,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd2,3'd1,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd4,3'd0,3'd1,3'd4,3'd0}};

parameter bit [2:0] SpriteTableG_3_14[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd4,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1},
'{3'd2,3'd2,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_3_15[7:0][7:0] = '{'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3},
'{3'd0,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd0,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd2,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3}};

parameter bit [2:0] SpriteTableG_3_16[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_3_17[7:0][7:0] = '{'{3'd3,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd3}};

parameter bit [2:0] SpriteTableG_3_18[7:0][7:0] = '{'{3'd1,3'd0,3'd0,3'd1,3'd2,3'd3,3'd3,3'd3},
'{3'd0,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_3_19[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd1,3'd2,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd0,3'd1,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_3_20[7:0][7:0] = '{'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd1,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_3_21[7:0][7:0] = '{'{3'd3,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_3_22[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd0,3'd2,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_3_23[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2},
'{3'd3,3'd3,3'd3,3'd2,3'd1,3'd0,3'd0,3'd0},
'{3'd2,3'd1,3'd0,3'd0,3'd1,3'd2,3'd2,3'd1},
'{3'd1,3'd1,3'd1,3'd0,3'd1,3'd3,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_3_24[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0},
'{3'd1,3'd3,3'd0,3'd0,3'd1,3'd3,3'd1,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd4,3'd3,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd0,3'd0,3'd2,3'd3,3'd2,3'd1},
'{3'd4,3'd1,3'd0,3'd1,3'd1,3'd3,3'd2,3'd1}};

parameter bit [2:0] SpriteTableG_3_25[7:0][7:0] = '{'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd4,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd2},
'{3'd2,3'd3,3'd2,3'd2,3'd2,3'd3,3'd3,3'd2},
'{3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd0,3'd2,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd0,3'd1,3'd3,3'd3,3'd2,3'd2,3'd2,3'd3},
'{3'd0,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_3_26[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd4,3'd1,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd1,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd1}};

parameter bit [2:0] SpriteTableG_3_27[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd3,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd3,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3},
'{3'd3,3'd3,3'd0,3'd0,3'd0,3'd0,3'd3,3'd3},
'{3'd3,3'd3,3'd4,3'd0,3'd0,3'd1,3'd3,3'd4},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd1,3'd1,3'd0}};

parameter bit [2:0] SpriteTableG_3_28[7:0][7:0] = '{'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd4,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd2,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_3_29[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd1,3'd1,3'd4,3'd4,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_3_30[7:0][7:0] = '{'{3'd0,3'd4,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd1},
'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1}};

parameter bit [2:0] SpriteTableG_3_31[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd1}};

parameter bit [2:0] SpriteTableG_3_32[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd3,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0},
'{3'd3,3'd3,3'd1,3'd3,3'd3,3'd4,3'd1,3'd2},
'{3'd4,3'd1,3'd3,3'd1,3'd0,3'd4,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4}};

parameter bit [2:0] SpriteTableG_3_33[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_3_34[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_3_35[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_4_0[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_4_1[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_4_2[7:0][7:0] = '{'{3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_4_3[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd2,3'd3,3'd3,3'd0},
'{3'd1,3'd0,3'd4,3'd2,3'd3,3'd3,3'd3,3'd0}};

parameter bit [2:0] SpriteTableG_4_4[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd3,3'd1,3'd1,3'd1}};

parameter bit [2:0] SpriteTableG_4_5[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd4,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd4,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd4,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd4,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd4,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_4_6[7:0][7:0] = '{'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd4,3'd3,3'd3,3'd1,3'd3},
'{3'd0,3'd0,3'd0,3'd4,3'd3,3'd2,3'd2,3'd2},
'{3'd0,3'd0,3'd4,3'd3,3'd2,3'd1,3'd1,3'd1},
'{3'd0,3'd1,3'd3,3'd3,3'd1,3'd1,3'd0,3'd1}};

parameter bit [2:0] SpriteTableG_4_7[7:0][7:0] = '{'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_4_8[7:0][7:0] = '{'{3'd3,3'd3,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd4,3'd0,3'd0,3'd0,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd2,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd1,3'd3,3'd3},
'{3'd1,3'd2,3'd3,3'd2,3'd1,3'd3,3'd3,3'd3},
'{3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_4_9[7:0][7:0] = '{'{3'd0,3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd2,3'd2,3'd3,3'd3},
'{3'd0,3'd1,3'd1,3'd4,3'd0,3'd0,3'd2,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_4_10[7:0][7:0] = '{'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd4,3'd2},
'{3'd0,3'd1,3'd1,3'd1,3'd2,3'd1,3'd2,3'd3},
'{3'd0,3'd0,3'd1,3'd1,3'd2,3'd2,3'd2,3'd3},
'{3'd0,3'd0,3'd1,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd1,3'd2,3'd3,3'd3,3'd2}};

parameter bit [2:0] SpriteTableG_4_11[7:0][7:0] = '{'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd2,3'd2,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd4,3'd0,3'd4,3'd2,3'd1}};

parameter bit [2:0] SpriteTableG_4_12[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_4_13[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd4,3'd3,3'd1},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd1,3'd3,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd1,3'd3,3'd0},
'{3'd0,3'd1,3'd3,3'd0,3'd0,3'd2,3'd1,3'd0}};

parameter bit [2:0] SpriteTableG_4_14[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1},
'{3'd0,3'd2,3'd3,3'd3,3'd3,3'd1,3'd3,3'd3},
'{3'd0,3'd0,3'd2,3'd3,3'd3,3'd1,3'd3,3'd3},
'{3'd0,3'd1,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_4_15[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3},
'{3'd0,3'd1,3'd1,3'd2,3'd2,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_4_16[7:0][7:0] = '{'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd0,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd1,3'd0,3'd2,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_4_17[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd3},
'{3'd0,3'd1,3'd0,3'd0,3'd0,3'd2,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0}};

parameter bit [2:0] SpriteTableG_4_18[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd1,3'd4,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_4_19[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_4_20[7:0][7:0] = '{'{3'd0,3'd0,3'd1,3'd0,3'd0,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd2,3'd3},
'{3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd1,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd1,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd2,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_4_21[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd0,3'd0,3'd2,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd0,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd0,3'd2,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd0,3'd2,3'd3,3'd3,3'd3,3'd3,3'd4,3'd0},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd1}};

parameter bit [2:0] SpriteTableG_4_22[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_4_23[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2},
'{3'd3,3'd3,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd3,3'd3,3'd1,3'd0,3'd2,3'd2,3'd2},
'{3'd0,3'd3,3'd3,3'd4,3'd0,3'd1,3'd3,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_4_24[7:0][7:0] = '{'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd4,3'd1,3'd1},
'{3'd4,3'd3,3'd3,3'd4,3'd0,3'd1,3'd3,3'd3},
'{3'd0,3'd3,3'd3,3'd4,3'd0,3'd1,3'd3,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd4,3'd4,3'd0,3'd0,3'd0,3'd1,3'd4},
'{3'd0,3'd3,3'd3,3'd0,3'd0,3'd1,3'd3,3'd1},
'{3'd0,3'd2,3'd1,3'd0,3'd0,3'd1,3'd3,3'd1}};

parameter bit [2:0] SpriteTableG_4_25[7:0][7:0] = '{'{3'd2,3'd3,3'd4,3'd0,3'd0,3'd0,3'd4,3'd4},
'{3'd2,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd3,3'd2,3'd0,3'd0,3'd0,3'd4,3'd0},
'{3'd2,3'd3,3'd3,3'd0,3'd0,3'd1,3'd3,3'd2},
'{3'd2,3'd3,3'd3,3'd0,3'd0,3'd2,3'd3,3'd2},
'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd1,3'd2,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd1,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd1}};

parameter bit [2:0] SpriteTableG_4_26[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd1,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd1,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd1,3'd1,3'd2},
'{3'd3,3'd3,3'd3,3'd1,3'd1,3'd0,3'd1,3'd1},
'{3'd3,3'd3,3'd2,3'd0,3'd0,3'd1,3'd3,3'd0},
'{3'd3,3'd3,3'd3,3'd0,3'd1,3'd3,3'd3,3'd4},
'{3'd3,3'd3,3'd2,3'd1,3'd3,3'd4,3'd1,3'd1}};

parameter bit [2:0] SpriteTableG_4_27[7:0][7:0] = '{'{3'd1,3'd3,3'd3,3'd3,3'd4,3'd0,3'd1,3'd1},
'{3'd0,3'd2,3'd3,3'd1,3'd0,3'd0,3'd0,3'd1},
'{3'd4,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_4_28[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd2},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1}};

parameter bit [2:0] SpriteTableG_4_29[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2},
'{3'd0,3'd0,3'd0,3'd4,3'd2,3'd2,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd4,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_4_30[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_4_31[7:0][7:0] = '{'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_4_32[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd3,3'd2,3'd1,3'd2,3'd4,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_4_33[7:0][7:0] = '{'{3'd3,3'd2,3'd1,3'd2,3'd2,3'd0,3'd0,3'd0},
'{3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_4_34[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_4_35[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_5_0[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_5_1[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_5_2[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1}};

parameter bit [2:0] SpriteTableG_5_3[7:0][7:0] = '{'{3'd0,3'd0,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_5_4[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd1,3'd4,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd4,3'd3,3'd3,3'd3},
'{3'd3,3'd2,3'd0,3'd0,3'd0,3'd2,3'd3,3'd3},
'{3'd3,3'd3,3'd2,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd3,3'd3,3'd2,3'd4,3'd0,3'd0,3'd2,3'd3}};

parameter bit [2:0] SpriteTableG_5_5[7:0][7:0] = '{'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd1,3'd0,3'd1,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd1,3'd4,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd4,3'd2,3'd3,3'd2,3'd2},
'{3'd0,3'd0,3'd0,3'd4,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd4,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd4,3'd1,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_5_6[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd1,3'd4,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd2,3'd1,3'd1,3'd0,3'd0},
'{3'd4,3'd1,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd3,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1}};

parameter bit [2:0] SpriteTableG_5_7[7:0][7:0] = '{'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_5_8[7:0][7:0] = '{'{3'd4,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd3,3'd2,3'd1,3'd2,3'd1,3'd0,3'd0},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_5_9[7:0][7:0] = '{'{3'd3,3'd3,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1}};

parameter bit [2:0] SpriteTableG_5_10[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd2},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd2},
'{3'd1,3'd0,3'd4,3'd4,3'd0,3'd0,3'd0,3'd1},
'{3'd1,3'd0,3'd1,3'd1,3'd0,3'd0,3'd4,3'd3},
'{3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_5_11[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd4,3'd1},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd1,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0},
'{3'd1,3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd0}};

parameter bit [2:0] SpriteTableG_5_12[7:0][7:0] = '{'{3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0},
'{3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0},
'{3'd1,3'd0,3'd1,3'd1,3'd0,3'd1,3'd0,3'd0},
'{3'd1,3'd0,3'd1,3'd0,3'd0,3'd1,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd1,3'd0,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd0,3'd1,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_5_13[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd0,3'd0,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd0,3'd0,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_5_14[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0},
'{3'd2,3'd2,3'd2,3'd2,3'd3,3'd2,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0},
'{3'd3,3'd3,3'd1,3'd1,3'd1,3'd4,3'd0,3'd0},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_5_15[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_5_16[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_5_17[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_5_18[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd4,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_5_19[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_5_20[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_5_21[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd4,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd1,3'd3},
'{3'd0,3'd4,3'd1,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_5_22[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd0}};

parameter bit [2:0] SpriteTableG_5_23[7:0][7:0] = '{'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd1,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0},
'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd1,3'd0},
'{3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd1,3'd0},
'{3'd0,3'd0,3'd1,3'd0,3'd1,3'd0,3'd1,3'd0},
'{3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd1,3'd0}};

parameter bit [2:0] SpriteTableG_5_24[7:0][7:0] = '{'{3'd1,3'd1,3'd2,3'd0,3'd1,3'd0,3'd1,3'd0},
'{3'd2,3'd2,3'd3,3'd0,3'd1,3'd0,3'd1,3'd0},
'{3'd1,3'd2,3'd3,3'd0,3'd1,3'd0,3'd1,3'd0},
'{3'd0,3'd2,3'd2,3'd0,3'd1,3'd0,3'd1,3'd0},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd0},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd0},
'{3'd0,3'd2,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1}};

parameter bit [2:0] SpriteTableG_5_25[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2},
'{3'd1,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd3},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd3},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd1,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1}};

parameter bit [2:0] SpriteTableG_5_26[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd3},
'{3'd0,3'd0,3'd1,3'd2,3'd1,3'd0,3'd1,3'd3},
'{3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd4,3'd1},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd2,3'd1,3'd0,3'd0,3'd4,3'd1},
'{3'd0,3'd1,3'd3,3'd3,3'd0,3'd0,3'd1,3'd3},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1}};

parameter bit [2:0] SpriteTableG_5_27[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd3},
'{3'd2,3'd1,3'd2,3'd2,3'd0,3'd0,3'd1,3'd3},
'{3'd2,3'd1,3'd1,3'd1,3'd2,3'd2,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd2,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2},
'{3'd0,3'd1,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_5_28[7:0][7:0] = '{'{3'd1,3'd2,3'd2,3'd0,3'd0,3'd2,3'd3,3'd3},
'{3'd1,3'd2,3'd3,3'd2,3'd1,3'd3,3'd1,3'd4},
'{3'd2,3'd1,3'd3,3'd3,3'd2,3'd1,3'd0,3'd0},
'{3'd2,3'd2,3'd2,3'd3,3'd2,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0},
'{3'd1,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd0},
'{3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd1,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_5_29[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd1,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_5_30[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4}};

parameter bit [2:0] SpriteTableG_5_31[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_5_32[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_5_33[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_5_34[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_5_35[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_6_0[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd3,3'd2,3'd1,3'd1,3'd4,3'd0}};

parameter bit [2:0] SpriteTableG_6_1[7:0][7:0] = '{'{3'd0,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd2,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_6_2[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd3,3'd3},
'{3'd1,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3},
'{3'd1,3'd0,3'd0,3'd0,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_6_3[7:0][7:0] = '{'{3'd1,3'd0,3'd0,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd0,3'd2,3'd3,3'd3,3'd3,3'd2,3'd2},
'{3'd0,3'd0,3'd2,3'd2,3'd1,3'd4,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd1,3'd2,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1}};

parameter bit [2:0] SpriteTableG_6_4[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd2,3'd3,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd2,3'd3,3'd3,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd3,3'd3,3'd3,3'd4,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1}};

parameter bit [2:0] SpriteTableG_6_5[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd0,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd1,3'd0,3'd1},
'{3'd2,3'd3,3'd3,3'd2,3'd1,3'd1,3'd0,3'd1},
'{3'd0,3'd1,3'd3,3'd2,3'd1,3'd1,3'd1,3'd2},
'{3'd0,3'd0,3'd2,3'd2,3'd1,3'd1,3'd1,3'd2},
'{3'd0,3'd0,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd1,3'd2,3'd1,3'd1,3'd1,3'd0,3'd4}};

parameter bit [2:0] SpriteTableG_6_6[7:0][7:0] = '{'{3'd0,3'd1,3'd4,3'd0,3'd1,3'd1,3'd2,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3},
'{3'd0,3'd0,3'd1,3'd1,3'd0,3'd4,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_6_7[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd3,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd3,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd3,3'd3,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd3,3'd3,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd3,3'd3,3'd0},
'{3'd1,3'd2,3'd1,3'd0,3'd4,3'd3,3'd3,3'd4},
'{3'd0,3'd2,3'd1,3'd0,3'd4,3'd3,3'd3,3'd4},
'{3'd0,3'd1,3'd4,3'd0,3'd0,3'd3,3'd3,3'd1}};

parameter bit [2:0] SpriteTableG_6_8[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd3,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd4,3'd3},
'{3'd0,3'd0,3'd0,3'd4,3'd1,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_6_9[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd2,3'd3,3'd1,3'd0,3'd0},
'{3'd4,3'd0,3'd0,3'd2,3'd3,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd2,3'd3,3'd1,3'd0,3'd0,3'd4},
'{3'd0,3'd0,3'd2,3'd3,3'd0,3'd0,3'd0,3'd1},
'{3'd4,3'd0,3'd3,3'd2,3'd0,3'd0,3'd4,3'd3}};

parameter bit [2:0] SpriteTableG_6_10[7:0][7:0] = '{'{3'd4,3'd0,3'd3,3'd1,3'd0,3'd0,3'd1,3'd3},
'{3'd4,3'd2,3'd2,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd1,3'd3,3'd2},
'{3'd3,3'd2,3'd0,3'd0,3'd0,3'd3,3'd3,3'd2},
'{3'd1,3'd1,3'd0,3'd0,3'd4,3'd3,3'd2,3'd2},
'{3'd4,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd2},
'{3'd0,3'd0,3'd0,3'd4,3'd3,3'd3,3'd3,3'd2},
'{3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd2}};

parameter bit [2:0] SpriteTableG_6_11[7:0][7:0] = '{'{3'd0,3'd4,3'd1,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd0,3'd0,3'd1,3'd3,3'd2,3'd2,3'd2,3'd2},
'{3'd0,3'd0,3'd1,3'd3,3'd2,3'd2,3'd3,3'd2},
'{3'd0,3'd0,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3},
'{3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd2,3'd2,3'd3,3'd2,3'd2},
'{3'd0,3'd1,3'd3,3'd3,3'd2,3'd3,3'd3,3'd2}};

parameter bit [2:0] SpriteTableG_6_12[7:0][7:0] = '{'{3'd0,3'd1,3'd3,3'd2,3'd2,3'd3,3'd3,3'd2},
'{3'd0,3'd3,3'd3,3'd2,3'd3,3'd2,3'd2,3'd2},
'{3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_6_13[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_6_14[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_6_15[7:0][7:0] = '{'{3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd4,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd0,3'd4,3'd1,3'd3,3'd3,3'd2,3'd3}};

parameter bit [2:0] SpriteTableG_6_16[7:0][7:0] = '{'{3'd3,3'd0,3'd0,3'd4,3'd3,3'd3,3'd0,3'd2},
'{3'd3,3'd4,3'd0,3'd0,3'd1,3'd3,3'd4,3'd0},
'{3'd3,3'd3,3'd0,3'd0,3'd4,3'd3,3'd3,3'd0},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd4,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd0,3'd0,3'd0,3'd4,3'd3},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd3,3'd3,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_6_17[7:0][7:0] = '{'{3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_6_18[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_6_19[7:0][7:0] = '{'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd4,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_6_20[7:0][7:0] = '{'{3'd3,3'd3,3'd4,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd1,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_6_21[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd3,3'd3,3'd3,3'd2},
'{3'd0,3'd0,3'd0,3'd4,3'd3,3'd3,3'd2,3'd3},
'{3'd1,3'd0,3'd0,3'd1,3'd3,3'd3,3'd2,3'd3},
'{3'd1,3'd0,3'd4,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd4,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_6_22[7:0][7:0] = '{'{3'd0,3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_6_23[7:0][7:0] = '{'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_6_24[7:0][7:0] = '{'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd4,3'd1,3'd3,3'd2,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_6_25[7:0][7:0] = '{'{3'd0,3'd0,3'd4,3'd3,3'd3,3'd2,3'd3,3'd3},
'{3'd4,3'd0,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd4,3'd4,3'd0,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd0,3'd1,3'd1,3'd0,3'd4,3'd1,3'd3,3'd3},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1}};

parameter bit [2:0] SpriteTableG_6_26[7:0][7:0] = '{'{3'd1,3'd0,3'd0,3'd1,3'd4,3'd0,3'd0,3'd0},
'{3'd3,3'd0,3'd4,3'd3,3'd3,3'd4,3'd0,3'd0},
'{3'd4,3'd0,3'd0,3'd1,3'd1,3'd4,3'd0,3'd0},
'{3'd0,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd1,3'd3,3'd4,3'd0,3'd1},
'{3'd1,3'd0,3'd0,3'd3,3'd3,3'd4,3'd0,3'd1},
'{3'd4,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd4}};

parameter bit [2:0] SpriteTableG_6_27[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd4,3'd1,3'd0,3'd0,3'd0},
'{3'd2,3'd0,3'd0,3'd1,3'd3,3'd0,3'd0,3'd1},
'{3'd3,3'd3,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_6_28[7:0][7:0] = '{'{3'd3,3'd3,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd2,3'd4,3'd4,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_6_29[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1}};

parameter bit [2:0] SpriteTableG_6_30[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd2},
'{3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1}};

parameter bit [2:0] SpriteTableG_6_31[7:0][7:0] = '{'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_6_32[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_6_33[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_6_34[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_6_35[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_7_0[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_7_1[7:0][7:0] = '{'{3'd2,3'd2,3'd1,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_7_2[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_7_3[7:0][7:0] = '{'{3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd1,3'd1,3'd0,3'd1,3'd3,3'd3,3'd3},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd3},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd3},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_7_4[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd2,3'd2,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd2,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd2,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_7_5[7:0][7:0] = '{'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd4,3'd1,3'd3},
'{3'd1,3'd0,3'd0,3'd0,3'd1,3'd3,3'd1,3'd4}};

parameter bit [2:0] SpriteTableG_7_6[7:0][7:0] = '{'{3'd3,3'd4,3'd4,3'd3,3'd3,3'd4,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_7_7[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_7_8[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3},
'{3'd3,3'd1,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd3,3'd4,3'd0,3'd0,3'd4,3'd3,3'd3,3'd2},
'{3'd4,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd2}};

parameter bit [2:0] SpriteTableG_7_9[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd3,3'd3,3'd2,3'd2,3'd2},
'{3'd0,3'd0,3'd1,3'd3,3'd2,3'd2,3'd2,3'd2},
'{3'd4,3'd4,3'd3,3'd3,3'd2,3'd2,3'd3,3'd2},
'{3'd4,3'd3,3'd3,3'd3,3'd2,3'd2,3'd3,3'd2},
'{3'd1,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd3,3'd3,3'd2,3'd3,3'd2,3'd2,3'd2,3'd2},
'{3'd3,3'd2,3'd2,3'd3,3'd2,3'd2,3'd3,3'd2},
'{3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableG_7_10[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd3,3'd3,3'd2,3'd3,3'd3,3'd2},
'{3'd2,3'd2,3'd3,3'd3,3'd2,3'd2,3'd3,3'd2},
'{3'd2,3'd2,3'd3,3'd2,3'd2,3'd2,3'd2,3'd3},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3},
'{3'd2,3'd2,3'd2,3'd2,3'd3,3'd2,3'd3,3'd3},
'{3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_7_11[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3},
'{3'd2,3'd2,3'd3,3'd2,3'd2,3'd2,3'd3,3'd3},
'{3'd2,3'd2,3'd3,3'd2,3'd2,3'd2,3'd2,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3},
'{3'd3,3'd2,3'd3,3'd2,3'd2,3'd3,3'd2,3'd3},
'{3'd3,3'd2,3'd2,3'd3,3'd2,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_7_12[7:0][7:0] = '{'{3'd3,3'd2,3'd2,3'd3,3'd2,3'd3,3'd3,3'd3},
'{3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1}};

parameter bit [2:0] SpriteTableG_7_13[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0}};

parameter bit [2:0] SpriteTableG_7_14[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_7_15[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_7_16[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd4,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd1,3'd0,3'd0,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd4,3'd1,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_7_17[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_7_18[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd4,3'd0,3'd1,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_7_19[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_7_20[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_7_21[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_7_22[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1}};

parameter bit [2:0] SpriteTableG_7_23[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_7_24[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_7_25[7:0][7:0] = '{'{3'd2,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_7_26[7:0][7:0] = '{'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd4,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4},
'{3'd0,3'd4,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd0,3'd4,3'd4,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd1,3'd0,3'd1,3'd3,3'd1,3'd1,3'd1},
'{3'd3,3'd3,3'd0,3'd4,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd1,3'd0,3'd0,3'd1,3'd3,3'd1,3'd1}};

parameter bit [2:0] SpriteTableG_7_27[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd4,3'd0,3'd0,3'd1,3'd1,3'd4,3'd0},
'{3'd3,3'd1,3'd0,3'd0,3'd3,3'd3,3'd1,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd1,3'd3,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd1,3'd1}};

parameter bit [2:0] SpriteTableG_7_28[7:0][7:0] = '{'{3'd3,3'd1,3'd0,3'd1,3'd3,3'd3,3'd2,3'd1},
'{3'd1,3'd4,3'd0,3'd0,3'd2,3'd3,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd1},
'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_7_29[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd3},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd3,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd3,3'd1}};

parameter bit [2:0] SpriteTableG_7_30[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd3,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd3,3'd1,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd3,3'd3,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd3,3'd1,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd2,3'd3,3'd4,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd2,3'd3,3'd0,3'd0,3'd0},
'{3'd1,3'd2,3'd1,3'd3,3'd3,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd1,3'd3,3'd3,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_7_31[7:0][7:0] = '{'{3'd1,3'd2,3'd1,3'd3,3'd3,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd2,3'd2,3'd3,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd2,3'd2,3'd3,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd4,3'd2,3'd3,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd3,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4}};

parameter bit [2:0] SpriteTableG_7_32[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_7_33[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_7_34[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_7_35[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_8_0[7:0][7:0] = '{'{3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd3,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd2,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd2,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_8_1[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd2,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_8_2[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd3,3'd3,3'd2,3'd2,3'd3,3'd3,3'd2,3'd2}};

parameter bit [2:0] SpriteTableG_8_3[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd3},
'{3'd3,3'd3,3'd2,3'd3,3'd3,3'd1,3'd0,3'd0},
'{3'd3,3'd3,3'd2,3'd3,3'd2,3'd1,3'd1,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd1,3'd4,3'd4,3'd0,3'd0,3'd4,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_8_4[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_8_5[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4},
'{3'd0,3'd4,3'd1,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd1,3'd3,3'd3,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd1,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_8_6[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_8_7[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_8_8[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd2,3'd2},
'{3'd0,3'd4,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2},
'{3'd1,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd3,3'd2,3'd2,3'd2,3'd3,3'd2,3'd2,3'd3},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd3,3'd2,3'd2,3'd3,3'd2,3'd2,3'd3}};

parameter bit [2:0] SpriteTableG_8_9[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd3,3'd2,3'd2,3'd3,3'd2,3'd2,3'd3},
'{3'd2,3'd3,3'd2,3'd2,3'd3,3'd2,3'd2,3'd3},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3},
'{3'd2,3'd3,3'd2,3'd2,3'd3,3'd2,3'd3,3'd1},
'{3'd2,3'd3,3'd2,3'd2,3'd2,3'd3,3'd3,3'd4}};

parameter bit [2:0] SpriteTableG_8_10[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd1,3'd0},
'{3'd2,3'd3,3'd3,3'd2,3'd3,3'd3,3'd0,3'd0},
'{3'd2,3'd3,3'd2,3'd2,3'd3,3'd1,3'd0,3'd0},
'{3'd2,3'd2,3'd2,3'd3,3'd3,3'd0,3'd0,3'd0},
'{3'd2,3'd3,3'd2,3'd3,3'd1,3'd0,3'd0,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd3},
'{3'd3,3'd2,3'd3,3'd1,3'd0,3'd0,3'd4,3'd3},
'{3'd2,3'd3,3'd3,3'd1,3'd0,3'd0,3'd1,3'd3}};

parameter bit [2:0] SpriteTableG_8_11[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd0,3'd0,3'd0,3'd3,3'd3},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd3,3'd3,3'd0,3'd0,3'd0,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3},
'{3'd3,3'd1,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3},
'{3'd3,3'd4,3'd0,3'd0,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd4,3'd0,3'd4,3'd3,3'd3,3'd3,3'd1}};

parameter bit [2:0] SpriteTableG_8_12[7:0][7:0] = '{'{3'd1,3'd0,3'd0,3'd0,3'd4,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd0,3'd0,3'd4,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd0,3'd0,3'd4,3'd0,3'd1,3'd1,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_8_13[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd0,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_8_14[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd4,3'd1,3'd1,3'd1,3'd3,3'd3},
'{3'd0,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd4},
'{3'd0,3'd4,3'd4,3'd3,3'd3,3'd1,3'd0,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd4,3'd0,3'd0,3'd4,3'd0,3'd0,3'd4},
'{3'd3,3'd3,3'd4,3'd4,3'd1,3'd4,3'd1,3'd3}};

parameter bit [2:0] SpriteTableG_8_15[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_8_16[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd2,3'd1,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd0,3'd0,3'd0,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd4,3'd0}};

parameter bit [2:0] SpriteTableG_8_17[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd3,3'd1,3'd0,3'd0,3'd4,3'd4,3'd1,3'd3},
'{3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd3,3'd2},
'{3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd2,3'd2},
'{3'd0,3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd2}};

parameter bit [2:0] SpriteTableG_8_18[7:0][7:0] = '{'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd2,3'd3,3'd3,3'd2,3'd2,3'd3},
'{3'd0,3'd3,3'd2,3'd3,3'd3,3'd2,3'd2,3'd2},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_8_19[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_8_20[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd0,3'd1}};

parameter bit [2:0] SpriteTableG_8_21[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd1,3'd4,3'd0,3'd4,3'd3},
'{3'd3,3'd3,3'd3,3'd4,3'd0,3'd0,3'd1,3'd3},
'{3'd3,3'd3,3'd3,3'd0,3'd0,3'd4,3'd3,3'd3},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd3,3'd3,3'd4,3'd0,3'd0,3'd3,3'd3,3'd3},
'{3'd3,3'd1,3'd0,3'd0,3'd4,3'd3,3'd3,3'd3},
'{3'd3,3'd1,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3},
'{3'd3,3'd1,3'd0,3'd0,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_8_22[7:0][7:0] = '{'{3'd3,3'd0,3'd0,3'd4,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd4,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd0,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd1}};

parameter bit [2:0] SpriteTableG_8_23[7:0][7:0] = '{'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd0,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd0,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd4,3'd1,3'd3,3'd3,3'd3,3'd1,3'd4},
'{3'd0,3'd4,3'd0,3'd1,3'd1,3'd4,3'd0,3'd4},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd1,3'd0,3'd0,3'd4,3'd0,3'd4,3'd1}};

parameter bit [2:0] SpriteTableG_8_24[7:0][7:0] = '{'{3'd3,3'd3,3'd1,3'd1,3'd3,3'd1,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_8_25[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_8_26[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd1,3'd4,3'd0,3'd0,3'd0},
'{3'd4,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd1},
'{3'd0,3'd0,3'd0,3'd4,3'd1,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_8_27[7:0][7:0] = '{'{3'd0,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd1,3'd3,3'd1,3'd0,3'd0,3'd3,3'd3,3'd2},
'{3'd1,3'd3,3'd3,3'd0,3'd4,3'd3,3'd3,3'd2},
'{3'd1,3'd3,3'd1,3'd0,3'd0,3'd3,3'd3,3'd2},
'{3'd0,3'd4,3'd0,3'd0,3'd0,3'd4,3'd4,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd1,3'd4,3'd0,3'd0,3'd1,3'd1,3'd1}};

parameter bit [2:0] SpriteTableG_8_28[7:0][7:0] = '{'{3'd1,3'd3,3'd3,3'd0,3'd0,3'd3,3'd3,3'd2},
'{3'd1,3'd3,3'd1,3'd0,3'd0,3'd3,3'd3,3'd2},
'{3'd2,3'd1,3'd0,3'd0,3'd0,3'd4,3'd1,3'd2},
'{3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd4,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_8_29[7:0][7:0] = '{'{3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd4,3'd4,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd1,3'd1,3'd4,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_8_30[7:0][7:0] = '{'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_8_31[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd1,3'd0,3'd0},
'{3'd1,3'd1,3'd4,3'd1,3'd1,3'd4,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_8_32[7:0][7:0] = '{'{3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd4,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd1,3'd4,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd1,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_8_33[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_8_34[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_8_35[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_9_0[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0},
'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0}};

parameter bit [2:0] SpriteTableG_9_1[7:0][7:0] = '{'{3'd0,3'd0,3'd1,3'd2,3'd1,3'd1,3'd1,3'd0},
'{3'd0,3'd0,3'd4,3'd2,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd2,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd1,3'd2,3'd1,3'd1,3'd1,3'd0},
'{3'd0,3'd0,3'd2,3'd1,3'd1,3'd1,3'd1,3'd0},
'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0},
'{3'd3,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_9_2[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd4,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd1,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0}};

parameter bit [2:0] SpriteTableG_9_3[7:0][7:0] = '{'{3'd3,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0},
'{3'd3,3'd3,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd1,3'd3,3'd2,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd3,3'd1,3'd2,3'd4,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd4,3'd1,3'd3,3'd3,3'd1,3'd4,3'd0},
'{3'd0,3'd0,3'd0,3'd4,3'd3,3'd3,3'd1,3'd4}};

parameter bit [2:0] SpriteTableG_9_4[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd1,3'd3,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_9_5[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd4,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_9_6[7:0][7:0] = '{'{3'd0,3'd0,3'd4,3'd4,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd4,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd4,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd3,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1}};

parameter bit [2:0] SpriteTableG_9_7[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4},
'{3'd0,3'd0,3'd4,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableG_9_8[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd3,3'd2,3'd2,3'd3,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd3,3'd2,3'd2,3'd3,3'd2,3'd2}};

parameter bit [2:0] SpriteTableG_9_9[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd2,3'd3,3'd3,3'd3,3'd1,3'd1,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd0,3'd0,3'd0,3'd4,3'd3},
'{3'd3,3'd3,3'd4,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd3,3'd0,3'd0,3'd0,3'd4,3'd0,3'd0,3'd0},
'{3'd4,3'd0,3'd0,3'd4,3'd3,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd3,3'd3,3'd3,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd4,3'd0}};

parameter bit [2:0] SpriteTableG_9_10[7:0][7:0] = '{'{3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd2,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd0,3'd2,3'd3}};

parameter bit [2:0] SpriteTableG_9_11[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd0,3'd0,3'd2,3'd3},
'{3'd3,3'd3,3'd3,3'd2,3'd0,3'd0,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd3,3'd3,3'd2,3'd0,3'd0,3'd2,3'd3,3'd3},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_9_12[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_9_13[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd1,3'd1,3'd4,3'd4,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_9_14[7:0][7:0] = '{'{3'd4,3'd0,3'd4,3'd0,3'd1,3'd3,3'd3,3'd3},
'{3'd1,3'd0,3'd4,3'd0,3'd3,3'd3,3'd3,3'd1},
'{3'd4,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd2},
'{3'd0,3'd4,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_9_15[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_9_16[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd4,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4}};

parameter bit [2:0] SpriteTableG_9_17[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd3,3'd3},
'{3'd0,3'd4,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd4,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3},
'{3'd2,3'd2,3'd3,3'd3,3'd3,3'd2,3'd2,3'd3},
'{3'd3,3'd3,3'd3,3'd2,3'd2,3'd1,3'd1,3'd2},
'{3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3}};

parameter bit [2:0] SpriteTableG_9_18[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd3,3'd3,3'd2,3'd2,3'd3},
'{3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd2,3'd3},
'{3'd3,3'd3,3'd2,3'd3,3'd3,3'd2,3'd2,3'd3},
'{3'd3,3'd2,3'd2,3'd3,3'd3,3'd0,3'd1,3'd3},
'{3'd2,3'd2,3'd3,3'd3,3'd3,3'd2,3'd1,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_9_19[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd1},
'{3'd3,3'd3,3'd3,3'd1,3'd4,3'd4,3'd0,3'd0},
'{3'd3,3'd3,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_9_20[7:0][7:0] = '{'{3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd1},
'{3'd0,3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd0,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_9_21[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_9_22[7:0][7:0] = '{'{3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd4,3'd0,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_9_23[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd3,3'd3},
'{3'd0,3'd0,3'd4,3'd0,3'd4,3'd3,3'd3,3'd3},
'{3'd1,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3},
'{3'd4,3'd0,3'd0,3'd4,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd4,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_9_24[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_9_25[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd4,3'd0,3'd0,3'd0,3'd1},
'{3'd3,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd3},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_9_26[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd4,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd2,3'd0,3'd2,3'd3,3'd3},
'{3'd2,3'd1,3'd0,3'd0,3'd0,3'd2,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_9_27[7:0][7:0] = '{'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd2,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd1,3'd0,3'd2,3'd3,3'd3},
'{3'd0,3'd1,3'd0,3'd1,3'd0,3'd3,3'd3,3'd1},
'{3'd0,3'd1,3'd0,3'd0,3'd0,3'd2,3'd1,3'd0},
'{3'd0,3'd1,3'd0,3'd0,3'd1,3'd0,3'd0,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd2},
'{3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd4}};

parameter bit [2:0] SpriteTableG_9_28[7:0][7:0] = '{'{3'd0,3'd0,3'd1,3'd0,3'd1,3'd3,3'd3,3'd0},
'{3'd0,3'd1,3'd0,3'd1,3'd3,3'd3,3'd4,3'd0},
'{3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd0,3'd0},
'{3'd0,3'd0,3'd4,3'd1,3'd3,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd3,3'd4,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3}};

parameter bit [2:0] SpriteTableG_9_29[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_9_30[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_9_31[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd4,3'd0}};

parameter bit [2:0] SpriteTableG_9_32[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd1},
'{3'd0,3'd0,3'd0,3'd4,3'd4,3'd1,3'd2,3'd4},
'{3'd4,3'd4,3'd4,3'd4,3'd1,3'd2,3'd2,3'd1},
'{3'd2,3'd1,3'd1,3'd1,3'd2,3'd3,3'd2,3'd1}};

parameter bit [2:0] SpriteTableG_9_33[7:0][7:0] = '{'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2},
'{3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd1,3'd3,3'd3,3'd2,3'd2,3'd3,3'd3,3'd2},
'{3'd1,3'd2,3'd4,3'd0,3'd0,3'd2,3'd3,3'd2}};

parameter bit [2:0] SpriteTableG_9_34[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_9_35[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_10_0[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_10_1[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3}};

parameter bit [2:0] SpriteTableG_10_2[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd3},
'{3'd0,3'd0,3'd0,3'd4,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd3,3'd2,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_10_3[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_10_4[7:0][7:0] = '{'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd1,3'd0,3'd1,3'd1,3'd0,3'd0},
'{3'd1,3'd3,3'd3,3'd0,3'd1,3'd1,3'd1,3'd0},
'{3'd4,3'd3,3'd3,3'd4,3'd1,3'd1,3'd1,3'd0},
'{3'd0,3'd1,3'd3,3'd1,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableG_10_5[7:0][7:0] = '{'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd3,3'd3,3'd3,3'd3,3'd1,3'd1,3'd1},
'{3'd3,3'd3,3'd1,3'd4,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_10_6[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_10_7[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd4,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd1,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3}};

parameter bit [2:0] SpriteTableG_10_8[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd3,3'd2,3'd2,3'd3,3'd2,3'd2,3'd3,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd3,3'd2,3'd2,3'd3,3'd2,3'd2,3'd3,3'd2}};

parameter bit [2:0] SpriteTableG_10_9[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd3,3'd2,3'd2,3'd3,3'd2,3'd2,3'd3,3'd2},
'{3'd3,3'd3,3'd2,3'd3,3'd2,3'd2,3'd3,3'd2},
'{3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd1,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd1}};

parameter bit [2:0] SpriteTableG_10_10[7:0][7:0] = '{'{3'd0,3'd1,3'd1,3'd1,3'd4,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4},
'{3'd0,3'd0,3'd4,3'd1,3'd1,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_10_11[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd1,3'd1,3'd4,3'd0,3'd0},
'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd0,3'd0,3'd1,3'd4,3'd0,3'd1,3'd4}};

parameter bit [2:0] SpriteTableG_10_12[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd4,3'd4,3'd1,3'd3,3'd3},
'{3'd1,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_10_13[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_10_14[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0}};

parameter bit [2:0] SpriteTableG_10_15[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd4,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd4,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd1,3'd1},
'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd1},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd4,3'd3},
'{3'd3,3'd3,3'd0,3'd0,3'd0,3'd4,3'd1,3'd3},
'{3'd3,3'd4,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3}};

parameter bit [2:0] SpriteTableG_10_16[7:0][7:0] = '{'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd0,3'd3,3'd1,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd4,3'd1,3'd4,3'd0,3'd0,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd4,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_10_17[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd3,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd2}};

parameter bit [2:0] SpriteTableG_10_18[7:0][7:0] = '{'{3'd3,3'd3,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd2,3'd2,3'd3,3'd3,3'd2},
'{3'd2,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_10_19[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_10_20[7:0][7:0] = '{'{3'd0,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd3,3'd2,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_10_21[7:0][7:0] = '{'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd2,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd1,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_10_22[7:0][7:0] = '{'{3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_10_23[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0}};

parameter bit [2:0] SpriteTableG_10_24[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd0,3'd1},
'{3'd3,3'd3,3'd3,3'd4,3'd0,3'd0,3'd1,3'd3},
'{3'd3,3'd3,3'd4,3'd0,3'd0,3'd4,3'd3,3'd3},
'{3'd3,3'd1,3'd0,3'd0,3'd0,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_10_25[7:0][7:0] = '{'{3'd1,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_10_26[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd1,3'd4,3'd0,3'd0,3'd4},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd1},
'{3'd3,3'd3,3'd3,3'd0,3'd0,3'd0,3'd4,3'd1},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd4,3'd1}};

parameter bit [2:0] SpriteTableG_10_27[7:0][7:0] = '{'{3'd3,3'd3,3'd4,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd2,3'd2,3'd0,3'd0,3'd0,3'd4,3'd1,3'd1},
'{3'd2,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1},
'{3'd2,3'd0,3'd0,3'd0,3'd0,3'd1,3'd4,3'd1},
'{3'd1,3'd0,3'd0,3'd0,3'd4,3'd1,3'd1,3'd1},
'{3'd4,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd4,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd4,3'd1,3'd4,3'd1,3'd1}};

parameter bit [2:0] SpriteTableG_10_28[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd1,3'd4,3'd1,3'd1,3'd4},
'{3'd0,3'd0,3'd4,3'd1,3'd4,3'd1,3'd1,3'd0},
'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0},
'{3'd0,3'd0,3'd1,3'd0,3'd1,3'd1,3'd1,3'd0},
'{3'd0,3'd4,3'd1,3'd0,3'd3,3'd1,3'd1,3'd0},
'{3'd0,3'd1,3'd1,3'd4,3'd1,3'd1,3'd4,3'd4},
'{3'd4,3'd1,3'd4,3'd1,3'd1,3'd1,3'd0,3'd1}};

parameter bit [2:0] SpriteTableG_10_29[7:0][7:0] = '{'{3'd3,3'd1,3'd0,3'd1,3'd1,3'd1,3'd0,3'd1},
'{3'd3,3'd1,3'd1,3'd3,3'd3,3'd3,3'd1,3'd3},
'{3'd3,3'd3,3'd3,3'd1,3'd1,3'd3,3'd3,3'd3},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_10_30[7:0][7:0] = '{'{3'd1,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_10_31[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_10_32[7:0][7:0] = '{'{3'd1,3'd4,3'd0,3'd0,3'd0,3'd4,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_10_33[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd4,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_10_34[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_10_35[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_11_0[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd2,3'd1,3'd1,3'd3,3'd1,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd4,3'd0},
'{3'd2,3'd2,3'd3,3'd3,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd3,3'd2,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_11_1[7:0][7:0] = '{'{3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0},
'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2}};

parameter bit [2:0] SpriteTableG_11_2[7:0][7:0] = '{'{3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd2},
'{3'd3,3'd3,3'd2,3'd4,3'd0,3'd0,3'd0,3'd1},
'{3'd3,3'd3,3'd3,3'd4,3'd0,3'd0,3'd0,3'd1},
'{3'd3,3'd2,3'd0,3'd0,3'd0,3'd0,3'd4,3'd2},
'{3'd3,3'd2,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2},
'{3'd3,3'd2,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd1,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_11_3[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3}};

parameter bit [2:0] SpriteTableG_11_4[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd3,3'd3},
'{3'd0,3'd4,3'd1,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd2,3'd3,3'd2,3'd2,3'd2,3'd2,3'd3}};

parameter bit [2:0] SpriteTableG_11_5[7:0][7:0] = '{'{3'd3,3'd3,3'd2,3'd1,3'd1,3'd2,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd2,3'd3,3'd3},
'{3'd0,3'd4,3'd1,3'd3,3'd3,3'd1,3'd1,3'd2},
'{3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd1,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd2,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3}};

parameter bit [2:0] SpriteTableG_11_6[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1}};

parameter bit [2:0] SpriteTableG_11_7[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd3,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd0,3'd0},
'{3'd0,3'd0,3'd4,3'd1,3'd3,3'd3,3'd4,3'd0},
'{3'd0,3'd0,3'd4,3'd3,3'd3,3'd3,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd3,3'd3,3'd1,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd4,3'd3,3'd3,3'd1},
'{3'd3,3'd1,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_11_8[7:0][7:0] = '{'{3'd2,3'd3,3'd1,3'd0,3'd0,3'd0,3'd3,3'd3},
'{3'd2,3'd3,3'd3,3'd1,3'd0,3'd0,3'd4,3'd3},
'{3'd2,3'd2,3'd3,3'd3,3'd0,3'd0,3'd0,3'd3},
'{3'd2,3'd2,3'd2,3'd3,3'd1,3'd0,3'd0,3'd1},
'{3'd2,3'd3,3'd2,3'd3,3'd3,3'd0,3'd0,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd3,3'd4,3'd0,3'd0},
'{3'd2,3'd2,3'd2,3'd2,3'd3,3'd1,3'd0,3'd0},
'{3'd2,3'd3,3'd2,3'd2,3'd3,3'd3,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_11_9[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd0,3'd0},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd4,3'd0},
'{3'd2,3'd3,3'd2,3'd2,3'd3,3'd3,3'd4,3'd0},
'{3'd2,3'd3,3'd2,3'd2,3'd3,3'd3,3'd1,3'd0},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd1,3'd1,3'd4,3'd0,3'd0},
'{3'd1,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_11_10[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd4,3'd1,3'd1,3'd3,3'd1},
'{3'd1,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0},
'{3'd3,3'd3,3'd1,3'd3,3'd1,3'd1,3'd0,3'd0},
'{3'd4,3'd0,3'd0,3'd4,3'd1,3'd1,3'd4,3'd0},
'{3'd4,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_11_11[7:0][7:0] = '{'{3'd1,3'd0,3'd0,3'd0,3'd4,3'd1,3'd0,3'd4},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd4,3'd0,3'd0},
'{3'd0,3'd1,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd0,3'd0,3'd4,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd3}};

parameter bit [2:0] SpriteTableG_11_12[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd4,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd1,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd4,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd0,3'd1,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd0,3'd1,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd1,3'd1,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd1,3'd4,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_11_13[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd4,3'd4,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd4,3'd1,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd0,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd1,3'd0,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd1,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd1,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd1,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_11_14[7:0][7:0] = '{'{3'd3,3'd1,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_11_15[7:0][7:0] = '{'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_11_16[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd1,3'd1,3'd1,3'd1,3'd4},
'{3'd4,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd1,3'd1,3'd0}};

parameter bit [2:0] SpriteTableG_11_17[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd0},
'{3'd3,3'd4,3'd0,3'd0,3'd0,3'd1,3'd3,3'd0},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd4,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd4,3'd0,3'd0},
'{3'd2,3'd3,3'd3,3'd2,3'd3,3'd1,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_11_18[7:0][7:0] = '{'{3'd2,3'd3,3'd3,3'd2,3'd3,3'd3,3'd0,3'd0},
'{3'd2,3'd3,3'd2,3'd2,3'd3,3'd3,3'd1,3'd0},
'{3'd2,3'd3,3'd3,3'd2,3'd3,3'd3,3'd1,3'd0},
'{3'd2,3'd3,3'd3,3'd2,3'd2,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1}};

parameter bit [2:0] SpriteTableG_11_19[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3},
'{3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd1}};

parameter bit [2:0] SpriteTableG_11_20[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4}};

parameter bit [2:0] SpriteTableG_11_21[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd1}};

parameter bit [2:0] SpriteTableG_11_22[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd0,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd4},
'{3'd3,3'd3,3'd3,3'd4,3'd0,3'd0,3'd0,3'd1},
'{3'd3,3'd3,3'd3,3'd0,3'd0,3'd0,3'd0,3'd1}};

parameter bit [2:0] SpriteTableG_11_23[7:0][7:0] = '{'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd3},
'{3'd3,3'd3,3'd4,3'd0,3'd0,3'd0,3'd0,3'd3},
'{3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3},
'{3'd3,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3},
'{3'd1,3'd0,3'd0,3'd4,3'd4,3'd0,3'd4,3'd3},
'{3'd4,3'd4,3'd0,3'd1,3'd4,3'd0,3'd4,3'd3},
'{3'd0,3'd0,3'd4,3'd3,3'd4,3'd0,3'd4,3'd3},
'{3'd0,3'd0,3'd1,3'd3,3'd0,3'd0,3'd1,3'd3}};

parameter bit [2:0] SpriteTableG_11_24[7:0][7:0] = '{'{3'd0,3'd4,3'd3,3'd3,3'd0,3'd0,3'd1,3'd3},
'{3'd0,3'd3,3'd3,3'd3,3'd0,3'd0,3'd1,3'd3},
'{3'd1,3'd3,3'd3,3'd1,3'd0,3'd0,3'd1,3'd3},
'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd1,3'd3},
'{3'd3,3'd3,3'd3,3'd4,3'd0,3'd0,3'd1,3'd3},
'{3'd3,3'd3,3'd4,3'd0,3'd0,3'd0,3'd1,3'd3},
'{3'd3,3'd3,3'd4,3'd0,3'd0,3'd0,3'd3,3'd3},
'{3'd3,3'd3,3'd1,3'd0,3'd4,3'd0,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_11_25[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd4,3'd0,3'd0,3'd3,3'd3},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd4,3'd3,3'd2},
'{3'd3,3'd1,3'd0,3'd0,3'd4,3'd1,3'd3,3'd1},
'{3'd3,3'd0,3'd4,3'd0,3'd4,3'd1,3'd3,3'd3},
'{3'd4,3'd0,3'd4,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd0,3'd4,3'd4,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd0,3'd4,3'd4,3'd0,3'd1,3'd1,3'd3,3'd3},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd1,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_11_26[7:0][7:0] = '{'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd4,3'd1,3'd4,3'd0,3'd0,3'd3,3'd3,3'd3},
'{3'd1,3'd1,3'd4,3'd0,3'd0,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd1,3'd1,3'd0,3'd4,3'd1,3'd3,3'd2,3'd3},
'{3'd1,3'd1,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_11_27[7:0][7:0] = '{'{3'd1,3'd4,3'd0,3'd3,3'd2,3'd2,3'd3,3'd3},
'{3'd1,3'd4,3'd2,3'd2,3'd1,3'd2,3'd2,3'd2},
'{3'd1,3'd4,3'd2,3'd1,3'd3,3'd3,3'd2,3'd2},
'{3'd1,3'd4,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd0,3'd0,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd4,3'd1,3'd4,3'd4,3'd1,3'd1,3'd4,3'd1},
'{3'd0,3'd1,3'd4,3'd0,3'd4,3'd4,3'd0,3'd0},
'{3'd4,3'd1,3'd0,3'd1,3'd3,3'd3,3'd1,3'd4}};

parameter bit [2:0] SpriteTableG_11_28[7:0][7:0] = '{'{3'd4,3'd3,3'd0,3'd3,3'd3,3'd3,3'd1,3'd1},
'{3'd1,3'd3,3'd0,3'd1,3'd3,3'd3,3'd1,3'd4},
'{3'd1,3'd1,3'd0,3'd4,3'd1,3'd1,3'd0,3'd0},
'{3'd1,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd1,3'd0,3'd4,3'd3,3'd1,3'd4,3'd0},
'{3'd3,3'd3,3'd0,3'd1,3'd3,3'd3,3'd1,3'd4},
'{3'd3,3'd3,3'd1,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_11_29[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0},
'{3'd0,3'd0,3'd0,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd3,3'd3,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd3,3'd1,3'd0}};

parameter bit [2:0] SpriteTableG_11_30[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd3,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3}};

parameter bit [2:0] SpriteTableG_11_31[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd3,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd4,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd3,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd3,3'd1,3'd0,3'd0,3'd0},
'{3'd4,3'd1,3'd3,3'd1,3'd3,3'd1,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_11_32[7:0][7:0] = '{'{3'd3,3'd3,3'd1,3'd0,3'd1,3'd1,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4},
'{3'd0,3'd4,3'd0,3'd0,3'd4,3'd2,3'd2,3'd0},
'{3'd0,3'd1,3'd2,3'd1,3'd2,3'd3,3'd2,3'd0},
'{3'd0,3'd0,3'd2,3'd2,3'd3,3'd3,3'd2,3'd0},
'{3'd0,3'd0,3'd1,3'd2,3'd2,3'd3,3'd2,3'd2}};

parameter bit [2:0] SpriteTableG_11_33[7:0][7:0] = '{'{3'd0,3'd0,3'd2,3'd3,3'd2,3'd2,3'd2,3'd2},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd2,3'd4},
'{3'd0,3'd1,3'd2,3'd1,3'd3,3'd3,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd3,3'd4,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd4,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd0,3'd0,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_11_34[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_11_35[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_12_0[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_12_1[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0}};

parameter bit [2:0] SpriteTableG_12_2[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_12_3[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_12_4[7:0][7:0] = '{'{3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd4,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd3,3'd4},
'{3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd0},
'{3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd4,3'd0}};

parameter bit [2:0] SpriteTableG_12_5[7:0][7:0] = '{'{3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd0},
'{3'd2,3'd3,3'd2,3'd2,3'd2,3'd3,3'd2,3'd0},
'{3'd2,3'd3,3'd2,3'd2,3'd2,3'd3,3'd3,3'd1},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1}};

parameter bit [2:0] SpriteTableG_12_6[7:0][7:0] = '{'{3'd2,3'd3,3'd1,3'd1,3'd1,3'd3,3'd2,3'd1},
'{3'd2,3'd3,3'd2,3'd1,3'd1,3'd3,3'd3,3'd1},
'{3'd2,3'd2,3'd1,3'd1,3'd1,3'd2,3'd2,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0},
'{3'd2,3'd3,3'd2,3'd1,3'd1,3'd3,3'd3,3'd0},
'{3'd3,3'd3,3'd2,3'd1,3'd2,3'd3,3'd3,3'd4},
'{3'd4,3'd1,3'd1,3'd1,3'd1,3'd3,3'd2,3'd0}};

parameter bit [2:0] SpriteTableG_12_7[7:0][7:0] = '{'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd1,3'd3,3'd4,3'd0,3'd1,3'd3,3'd3,3'd0},
'{3'd3,3'd3,3'd3,3'd0,3'd1,3'd3,3'd3,3'd1},
'{3'd1,3'd3,3'd1,3'd0,3'd4,3'd1,3'd1,3'd0},
'{3'd0,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1}};

parameter bit [2:0] SpriteTableG_12_8[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd0,3'd0,3'd0,3'd0,3'd3},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd4,3'd3},
'{3'd3,3'd3,3'd3,3'd0,3'd0,3'd0,3'd1,3'd3},
'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd4,3'd0,3'd4,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd0,3'd0,3'd4,3'd3,3'd2},
'{3'd1,3'd3,3'd1,3'd0,3'd0,3'd1,3'd3,3'd2},
'{3'd1,3'd3,3'd1,3'd0,3'd0,3'd3,3'd3,3'd2}};

parameter bit [2:0] SpriteTableG_12_9[7:0][7:0] = '{'{3'd4,3'd3,3'd4,3'd0,3'd0,3'd3,3'd3,3'd2},
'{3'd4,3'd1,3'd0,3'd0,3'd1,3'd3,3'd2,3'd2},
'{3'd4,3'd1,3'd0,3'd0,3'd1,3'd3,3'd2,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd3,3'd3,3'd2,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd3,3'd3,3'd2,3'd2},
'{3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd2,3'd2},
'{3'd0,3'd0,3'd4,3'd1,3'd3,3'd3,3'd3,3'd2},
'{3'd0,3'd0,3'd0,3'd3,3'd3,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableG_12_10[7:0][7:0] = '{'{3'd0,3'd0,3'd4,3'd3,3'd3,3'd2,3'd2,3'd2},
'{3'd0,3'd0,3'd1,3'd3,3'd2,3'd3,3'd3,3'd2},
'{3'd0,3'd0,3'd1,3'd3,3'd2,3'd3,3'd3,3'd2},
'{3'd0,3'd0,3'd3,3'd3,3'd2,3'd2,3'd3,3'd3},
'{3'd0,3'd4,3'd3,3'd3,3'd2,3'd3,3'd3,3'd2},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_12_11[7:0][7:0] = '{'{3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_12_12[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_12_13[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_12_14[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_12_15[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0}};

parameter bit [2:0] SpriteTableG_12_16[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd4,3'd0},
'{3'd3,3'd3,3'd3,3'd1,3'd1,3'd4,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_12_17[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd4,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd2,3'd2,3'd3,3'd2,3'd2},
'{3'd0,3'd1,3'd3,3'd2,3'd1,3'd1,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_12_18[7:0][7:0] = '{'{3'd0,3'd1,3'd3,3'd2,3'd1,3'd1,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd2,3'd1,3'd2,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd2,3'd3,3'd2,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd2,3'd2,3'd3,3'd2,3'd3},
'{3'd0,3'd1,3'd3,3'd2,3'd3,3'd3,3'd2,3'd2},
'{3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_12_19[7:0][7:0] = '{'{3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd3,3'd3,3'd2,3'd1,3'd3,3'd3,3'd3},
'{3'd4,3'd3,3'd3,3'd3,3'd1,3'd2,3'd3,3'd3},
'{3'd0,3'd3,3'd3,3'd3,3'd2,3'd2,3'd3,3'd3},
'{3'd4,3'd3,3'd3,3'd3,3'd3,3'd1,3'd3,3'd3},
'{3'd4,3'd3,3'd3,3'd3,3'd3,3'd4,3'd2,3'd3},
'{3'd4,3'd3,3'd3,3'd3,3'd3,3'd1,3'd2,3'd3}};

parameter bit [2:0] SpriteTableG_12_20[7:0][7:0] = '{'{3'd4,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_12_21[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_12_22[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2},
'{3'd1,3'd2,3'd3,3'd3,3'd3,3'd2,3'd0,3'd4}};

parameter bit [2:0] SpriteTableG_12_23[7:0][7:0] = '{'{3'd1,3'd1,3'd3,3'd3,3'd3,3'd2,3'd1,3'd2},
'{3'd1,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd0,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd4,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd1,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd2,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_12_24[7:0][7:0] = '{'{3'd3,3'd3,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd4,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd1,3'd4,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd2,3'd0,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_12_25[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_12_26[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd4,3'd1,3'd4},
'{3'd1,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd0,3'd1,3'd1},
'{3'd1,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_12_27[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd2,3'd2,3'd1,3'd1,3'd0},
'{3'd2,3'd3,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd2,3'd3,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd1,3'd3,3'd3,3'd0,3'd1},
'{3'd2,3'd3,3'd2,3'd1,3'd2,3'd3,3'd1,3'd0},
'{3'd1,3'd2,3'd1,3'd1,3'd1,3'd2,3'd2,3'd0},
'{3'd3,3'd3,3'd3,3'd1,3'd2,3'd3,3'd3,3'd2}};

parameter bit [2:0] SpriteTableG_12_28[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd1,3'd3,3'd3,3'd3,3'd1},
'{3'd1,3'd3,3'd2,3'd0,3'd4,3'd3,3'd1,3'd4},
'{3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd3,3'd1,3'd0,3'd1,3'd3,3'd3,3'd4},
'{3'd3,3'd3,3'd3,3'd0,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd0,3'd1,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd1,3'd0,3'd4,3'd3,3'd3,3'd4}};

parameter bit [2:0] SpriteTableG_12_29[7:0][7:0] = '{'{3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd1,3'd4,3'd0,3'd4,3'd1,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd0,3'd1,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd0,3'd1,3'd3,3'd3,3'd1},
'{3'd1,3'd3,3'd4,3'd0,3'd4,3'd3,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0},
'{3'd3,3'd3,3'd1,3'd0,3'd1,3'd3,3'd3,3'd4}};

parameter bit [2:0] SpriteTableG_12_30[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd0,3'd1,3'd3,3'd3,3'd1},
'{3'd1,3'd3,3'd4,3'd0,3'd4,3'd3,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd0,3'd0},
'{3'd1,3'd3,3'd1,3'd0,3'd4,3'd3,3'd3,3'd4},
'{3'd3,3'd3,3'd1,3'd0,3'd1,3'd3,3'd3,3'd4},
'{3'd1,3'd3,3'd4,3'd0,3'd4,3'd3,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_12_31[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd4,3'd0,3'd0,3'd1,3'd1,3'd0},
'{3'd3,3'd3,3'd1,3'd0,3'd4,3'd3,3'd3,3'd4},
'{3'd1,3'd1,3'd4,3'd0,3'd0,3'd1,3'd3,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd3},
'{3'd0,3'd4,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd1,3'd3,3'd4,3'd0,3'd4,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_12_32[7:0][7:0] = '{'{3'd4,3'd1,3'd0,3'd0,3'd0,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd4,3'd1,3'd3,3'd3,3'd3,3'd2},
'{3'd2,3'd3,3'd2,3'd3,3'd3,3'd3,3'd2,3'd2},
'{3'd3,3'd3,3'd2,3'd2,3'd3,3'd2,3'd2,3'd3},
'{3'd1,3'd3,3'd3,3'd2,3'd2,3'd3,3'd3,3'd3},
'{3'd4,3'd1,3'd2,3'd3,3'd2,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd2,3'd3,3'd2,3'd2,3'd3},
'{3'd4,3'd4,3'd0,3'd4,3'd3,3'd3,3'd2,3'd2}};

parameter bit [2:0] SpriteTableG_12_33[7:0][7:0] = '{'{3'd1,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd2},
'{3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd2},
'{3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd2,3'd0},
'{3'd0,3'd0,3'd0,3'd2,3'd3,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd4,3'd0,3'd4,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd0,3'd0},
'{3'd4,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_12_34[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_12_35[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_13_0[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1}};

parameter bit [2:0] SpriteTableG_13_1[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd4,3'd0,3'd0,3'd0,3'd1,3'd3},
'{3'd0,3'd4,3'd3,3'd2,3'd2,3'd1,3'd3,3'd3},
'{3'd0,3'd0,3'd2,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_13_2[7:0][7:0] = '{'{3'd1,3'd0,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4},
'{3'd0,3'd4,3'd1,3'd0,3'd3,3'd3,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd3,3'd4,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd3,3'd3,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd4,3'd3,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd4,3'd3,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd3,3'd1,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_13_3[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd1,3'd3,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd4,3'd3,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd3,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd2,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_13_4[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_13_5[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd4,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd0,3'd4,3'd1,3'd4,3'd0,3'd0,3'd1,3'd2},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd1,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd1},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd4,3'd1,3'd0}};

parameter bit [2:0] SpriteTableG_13_6[7:0][7:0] = '{'{3'd1,3'd2,3'd3,3'd2,3'd1,3'd0,3'd1,3'd0},
'{3'd1,3'd2,3'd3,3'd1,3'd0,3'd4,3'd1,3'd0},
'{3'd1,3'd1,3'd4,3'd0,3'd0,3'd1,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0},
'{3'd0,3'd1,3'd3,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd3,3'd3,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd4,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_13_7[7:0][7:0] = '{'{3'd0,3'd1,3'd1,3'd2,3'd0,3'd0,3'd1,3'd0},
'{3'd0,3'd2,3'd3,3'd2,3'd0,3'd1,3'd0,3'd0},
'{3'd0,3'd1,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd3,3'd3,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd1},
'{3'd1,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_13_8[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd3,3'd2,3'd2,3'd3,3'd2,3'd2,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_13_9[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd3,3'd2,3'd2,3'd3,3'd2,3'd2,3'd3,3'd2},
'{3'd3,3'd3,3'd2,3'd3,3'd3,3'd2,3'd3,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3},
'{3'd3,3'd3,3'd2,3'd3,3'd3,3'd2,3'd3,3'd3},
'{3'd2,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3}};

parameter bit [2:0] SpriteTableG_13_10[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3},
'{3'd3,3'd3,3'd2,3'd3,3'd2,3'd2,3'd3,3'd3},
'{3'd3,3'd3,3'd2,3'd3,3'd3,3'd2,3'd3,3'd3},
'{3'd2,3'd2,3'd3,3'd3,3'd2,3'd2,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd1},
'{3'd3,3'd3,3'd2,3'd3,3'd2,3'd2,3'd3,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd3,3'd0}};

parameter bit [2:0] SpriteTableG_13_11[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd3,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd0}};

parameter bit [2:0] SpriteTableG_13_12[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd4,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd4,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd0,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd0,3'd0,3'd0,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd4,3'd1},
'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd1}};

parameter bit [2:0] SpriteTableG_13_13[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd4,3'd0,3'd0,3'd0,3'd1},
'{3'd3,3'd3,3'd3,3'd2,3'd1,3'd4,3'd1,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_13_14[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd1,3'd1,3'd1,3'd1,3'd1,3'd3,3'd3},
'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3},
'{3'd4,3'd4,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3}};

parameter bit [2:0] SpriteTableG_13_15[7:0][7:0] = '{'{3'd4,3'd4,3'd4,3'd4,3'd0,3'd0,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd3,3'd3},
'{3'd0,3'd0,3'd3,3'd1,3'd0,3'd0,3'd3,3'd3},
'{3'd0,3'd0,3'd3,3'd1,3'd0,3'd4,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd4,3'd0,3'd4,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd4,3'd0,3'd4,3'd3,3'd3},
'{3'd0,3'd3,3'd3,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd0,3'd3,3'd3,3'd0,3'd0,3'd1,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_13_16[7:0][7:0] = '{'{3'd4,3'd3,3'd3,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd1,3'd3,3'd1,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd1,3'd3,3'd1,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd4,3'd0,3'd0,3'd3,3'd3,3'd1},
'{3'd1,3'd4,3'd0,3'd0,3'd0,3'd0,3'd4,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_13_17[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_13_18[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd4},
'{3'd3,3'd4,3'd1,3'd3,3'd3,3'd3,3'd3,3'd4},
'{3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4}};

parameter bit [2:0] SpriteTableG_13_19[7:0][7:0] = '{'{3'd0,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd2,3'd3,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd2,3'd3,3'd3,3'd1,3'd0}};

parameter bit [2:0] SpriteTableG_13_20[7:0][7:0] = '{'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd1,3'd4},
'{3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd4,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_13_21[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd4,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd4,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd3},
'{3'd2,3'd2,3'd3,3'd3,3'd3,3'd0,3'd1,3'd3},
'{3'd2,3'd0,3'd2,3'd3,3'd3,3'd0,3'd1,3'd3}};

parameter bit [2:0] SpriteTableG_13_22[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd1,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd4,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd4,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd1,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd1,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_13_23[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_13_24[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd1,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_13_25[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_13_26[7:0][7:0] = '{'{3'd3,3'd3,3'd1,3'd1,3'd1,3'd4,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd0,3'd0,3'd4,3'd1,3'd1,3'd1,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_13_27[7:0][7:0] = '{'{3'd0,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd0,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd0,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd1,3'd0,3'd1,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd0,3'd0,3'd0,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_13_28[7:0][7:0] = '{'{3'd0,3'd1,3'd0,3'd0,3'd0,3'd2,3'd3,3'd3},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd3,3'd3},
'{3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd2,3'd3},
'{3'd0,3'd2,3'd0,3'd1,3'd0,3'd0,3'd1,3'd3},
'{3'd4,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd2},
'{3'd4,3'd3,3'd3,3'd0,3'd1,3'd0,3'd0,3'd1},
'{3'd0,3'd1,3'd3,3'd1,3'd1,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_13_29[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd1,3'd0},
'{3'd0,3'd2,3'd3,3'd2,3'd0,3'd0,3'd1,3'd0},
'{3'd0,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0},
'{3'd4,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd3,3'd2,3'd1,3'd1,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd0,3'd4,3'd2,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd0,3'd3,3'd3,3'd3,3'd0,3'd2,3'd2,3'd1}};

parameter bit [2:0] SpriteTableG_13_30[7:0][7:0] = '{'{3'd0,3'd3,3'd3,3'd3,3'd0,3'd1,3'd3,3'd0},
'{3'd0,3'd1,3'd3,3'd1,3'd0,3'd4,3'd3,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd4,3'd0,3'd0,3'd0,3'd4,3'd1},
'{3'd0,3'd1,3'd3,3'd1,3'd0,3'd4,3'd3,3'd3},
'{3'd0,3'd3,3'd3,3'd3,3'd0,3'd2,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd1,3'd0,3'd1,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1}};

parameter bit [2:0] SpriteTableG_13_31[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd1,3'd3,3'd1,3'd1,3'd1,3'd3,3'd3},
'{3'd0,3'd3,3'd3,3'd1,3'd0,3'd2,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd1,3'd0,3'd1,3'd3,3'd1},
'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd1,3'd1,3'd4,3'd0,3'd0,3'd1,3'd1},
'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_13_32[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd2,3'd1,3'd1,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd1,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd0,3'd1,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_13_33[7:0][7:0] = '{'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd4,3'd1},
'{3'd1,3'd2,3'd3,3'd3,3'd3,3'd1,3'd4,3'd1},
'{3'd0,3'd0,3'd0,3'd1,3'd3,3'd2,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd0,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd2,3'd3,3'd4,3'd1,3'd2},
'{3'd0,3'd0,3'd0,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd2,3'd3,3'd3,3'd3,3'd2}};

parameter bit [2:0] SpriteTableG_13_34[7:0][7:0] = '{'{3'd0,3'd4,3'd2,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd2,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd2,3'd3,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_13_35[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_14_0[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd3,3'd3},
'{3'd0,3'd0,3'd4,3'd3,3'd3,3'd1,3'd1,3'd1},
'{3'd0,3'd1,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd3,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_14_1[7:0][7:0] = '{'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd1,3'd1,3'd4,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_14_2[7:0][7:0] = '{'{3'd1,3'd4,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_14_3[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd1,3'd4,3'd4,3'd0,3'd0,3'd0},
'{3'd2,3'd3,3'd1,3'd4,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd3,3'd3,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd4,3'd1,3'd1,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_14_4[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_14_5[7:0][7:0] = '{'{3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1},
'{3'd1,3'd0,3'd1,3'd1,3'd4,3'd0,3'd0,3'd2},
'{3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd1,3'd2},
'{3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd2,3'd3},
'{3'd0,3'd0,3'd0,3'd1,3'd0,3'd4,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_14_6[7:0][7:0] = '{'{3'd0,3'd1,3'd0,3'd2,3'd4,3'd1,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd3,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd2,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd1,3'd0,3'd1,3'd1,3'd0,3'd0,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_14_7[7:0][7:0] = '{'{3'd1,3'd0,3'd2,3'd2,3'd0,3'd0,3'd2,3'd3},
'{3'd0,3'd0,3'd2,3'd3,3'd0,3'd0,3'd3,3'd3},
'{3'd0,3'd0,3'd3,3'd3,3'd1,3'd1,3'd2,3'd1},
'{3'd1,3'd1,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_14_8[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd3,3'd3,3'd2,3'd3,3'd3,3'd2,3'd3}};

parameter bit [2:0] SpriteTableG_14_9[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd3,3'd3,3'd3,3'd2,3'd2,3'd3,3'd2,3'd3},
'{3'd3,3'd3,3'd3,3'd2,3'd3,3'd3,3'd2,3'd3},
'{3'd3,3'd1,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd3,3'd1,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd3,3'd1,3'd3,3'd2,3'd3,3'd3,3'd2,3'd3},
'{3'd1,3'd1,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableG_14_10[7:0][7:0] = '{'{3'd1,3'd1,3'd3,3'd2,3'd2,3'd2,3'd3,3'd2},
'{3'd4,3'd1,3'd3,3'd2,3'd2,3'd3,3'd2,3'd3},
'{3'd0,3'd1,3'd3,3'd2,3'd3,3'd3,3'd2,3'd3},
'{3'd0,3'd1,3'd3,3'd2,3'd3,3'd2,3'd2,3'd2},
'{3'd0,3'd1,3'd2,3'd2,3'd2,3'd3,3'd2,3'd2},
'{3'd0,3'd3,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3},
'{3'd0,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd3},
'{3'd4,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd3}};

parameter bit [2:0] SpriteTableG_14_11[7:0][7:0] = '{'{3'd4,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd3},
'{3'd4,3'd3,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3},
'{3'd1,3'd3,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd2,3'd3,3'd2,3'd3},
'{3'd1,3'd3,3'd3,3'd2,3'd3,3'd3,3'd2,3'd3}};

parameter bit [2:0] SpriteTableG_14_12[7:0][7:0] = '{'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_14_13[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_14_14[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_14_15[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_14_16[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd1,3'd1,3'd4},
'{3'd1,3'd1,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_14_17[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_14_18[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd4,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_14_19[7:0][7:0] = '{'{3'd0,3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd4,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_14_20[7:0][7:0] = '{'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_14_21[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_14_22[7:0][7:0] = '{'{3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd1,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_14_23[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd2,3'd1},
'{3'd3,3'd3,3'd2,3'd2,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd1,3'd3,3'd3,3'd3,3'd2},
'{3'd3,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3}};

parameter bit [2:0] SpriteTableG_14_24[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4},
'{3'd3,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd0},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd0}};

parameter bit [2:0] SpriteTableG_14_25[7:0][7:0] = '{'{3'd3,3'd2,3'd3,3'd2,3'd3,3'd3,3'd4,3'd0},
'{3'd3,3'd3,3'd2,3'd2,3'd3,3'd1,3'd0,3'd0},
'{3'd3,3'd3,3'd2,3'd3,3'd3,3'd1,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd0},
'{3'd2,3'd2,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd4,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd4,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_14_26[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd0,3'd0},
'{3'd4,3'd1,3'd1,3'd1,3'd3,3'd3,3'd4,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0}};

parameter bit [2:0] SpriteTableG_14_27[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_14_28[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd3,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1}};

parameter bit [2:0] SpriteTableG_14_29[7:0][7:0] = '{'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd0},
'{3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd0,3'd2,3'd3,3'd3,3'd3,3'd3,3'd0,3'd0},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd0,3'd0},
'{3'd1,3'd0,3'd3,3'd3,3'd3,3'd2,3'd0,3'd0},
'{3'd0,3'd0,3'd2,3'd3,3'd3,3'd2,3'd0,3'd1},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd1,3'd0,3'd2}};

parameter bit [2:0] SpriteTableG_14_30[7:0][7:0] = '{'{3'd1,3'd1,3'd0,3'd3,3'd3,3'd0,3'd0,3'd2},
'{3'd0,3'd0,3'd0,3'd2,3'd3,3'd0,3'd0,3'd3},
'{3'd0,3'd1,3'd0,3'd1,3'd2,3'd0,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd1,3'd4},
'{3'd1,3'd0,3'd1,3'd0,3'd0,3'd0,3'd1,3'd3},
'{3'd2,3'd0,3'd0,3'd1,3'd1,3'd0,3'd2,3'd3},
'{3'd1,3'd0,3'd0,3'd1,3'd0,3'd0,3'd4,3'd3},
'{3'd0,3'd1,3'd0,3'd1,3'd0,3'd1,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_14_31[7:0][7:0] = '{'{3'd0,3'd1,3'd0,3'd1,3'd0,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd1,3'd1},
'{3'd1,3'd0,3'd1,3'd0,3'd0,3'd2,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd0,3'd1,3'd2,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd3,3'd3},
'{3'd0,3'd0,3'd4,3'd2,3'd1,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_14_32[7:0][7:0] = '{'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd4,3'd1,3'd1,3'd2,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd0,3'd0,3'd4,3'd3,3'd4,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd4,3'd3,3'd4,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_14_33[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_14_34[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_14_35[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_15_0[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd4,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd4,3'd3,3'd3,3'd4,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd3,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd3,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd3,3'd1,3'd4}};

parameter bit [2:0] SpriteTableG_15_1[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd1,3'd0,3'd0},
'{3'd0,3'd4,3'd1,3'd4,3'd1,3'd0,3'd0,3'd0},
'{3'd4,3'd4,3'd4,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd4,3'd0,3'd0,3'd0,3'd1,3'd4,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd4,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_15_2[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd4,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd4,3'd4,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_15_3[7:0][7:0] = '{'{3'd0,3'd0,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd4,3'd4,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd4,3'd1,3'd3,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd2,3'd1},
'{3'd0,3'd0,3'd0,3'd1,3'd3,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd3,3'd3,3'd2,3'd1,3'd1,3'd1},
'{3'd3,3'd3,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1}};

parameter bit [2:0] SpriteTableG_15_4[7:0][7:0] = '{'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd1},
'{3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_15_5[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd4,3'd3,3'd4,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd4,3'd3,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_15_6[7:0][7:0] = '{'{3'd3,3'd0,3'd0,3'd0,3'd4,3'd4,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd1,3'd3,3'd0,3'd4},
'{3'd3,3'd2,3'd1,3'd1,3'd2,3'd1,3'd0,3'd0},
'{3'd3,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd3,3'd3,3'd2,3'd1,3'd1,3'd0,3'd2,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd4,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd3}};

parameter bit [2:0] SpriteTableG_15_7[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd2,3'd2,3'd1,3'd1,3'd0},
'{3'd1,3'd4,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd2,3'd1},
'{3'd1,3'd1,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_15_8[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd1},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd1},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd1},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd1},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd1},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd1},
'{3'd3,3'd2,3'd3,3'd3,3'd2,3'd2,3'd3,3'd1}};

parameter bit [2:0] SpriteTableG_15_9[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd1},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd4},
'{3'd3,3'd2,3'd2,3'd3,3'd2,3'd3,3'd3,3'd4},
'{3'd3,3'd2,3'd3,3'd3,3'd2,3'd3,3'd3,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd0},
'{3'd3,3'd2,3'd3,3'd3,3'd2,3'd3,3'd3,3'd0},
'{3'd3,3'd2,3'd2,3'd3,3'd2,3'd3,3'd3,3'd0}};

parameter bit [2:0] SpriteTableG_15_10[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd0},
'{3'd2,3'd2,3'd3,3'd3,3'd2,3'd3,3'd3,3'd0},
'{3'd2,3'd2,3'd3,3'd3,3'd2,3'd3,3'd3,3'd0},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd1,3'd0},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd1,3'd0},
'{3'd2,3'd2,3'd3,3'd3,3'd2,3'd3,3'd1,3'd0},
'{3'd2,3'd2,3'd3,3'd3,3'd2,3'd3,3'd1,3'd0},
'{3'd2,3'd2,3'd3,3'd3,3'd2,3'd3,3'd1,3'd0}};

parameter bit [2:0] SpriteTableG_15_11[7:0][7:0] = '{'{3'd2,3'd2,3'd3,3'd3,3'd2,3'd3,3'd1,3'd0},
'{3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd1,3'd0},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd1,3'd0},
'{3'd3,3'd2,3'd2,3'd1,3'd2,3'd3,3'd1,3'd0}};

parameter bit [2:0] SpriteTableG_15_12[7:0][7:0] = '{'{3'd3,3'd2,3'd3,3'd2,3'd2,3'd3,3'd1,3'd0},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd0},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd0}};

parameter bit [2:0] SpriteTableG_15_13[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd1}};

parameter bit [2:0] SpriteTableG_15_14[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd1,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd1,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_15_15[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_15_16[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_15_17[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd4,3'd4,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_15_18[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_15_19[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd2,3'd2,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0}};

parameter bit [2:0] SpriteTableG_15_20[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd4,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd4}};

parameter bit [2:0] SpriteTableG_15_21[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd0,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd4,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd0,3'd0,3'd0,3'd3},
'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd3},
'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd1,3'd3},
'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd4,3'd1,3'd3}};

parameter bit [2:0] SpriteTableG_15_22[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd4,3'd0,3'd0,3'd1,3'd3},
'{3'd3,3'd3,3'd3,3'd0,3'd0,3'd0,3'd1,3'd3},
'{3'd3,3'd3,3'd3,3'd4,3'd0,3'd1,3'd3,3'd3},
'{3'd3,3'd3,3'd1,3'd4,3'd0,3'd4,3'd3,3'd3},
'{3'd3,3'd3,3'd4,3'd0,3'd0,3'd4,3'd3,3'd3},
'{3'd3,3'd3,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd3,3'd3,3'd0,3'd4,3'd0,3'd1,3'd3,3'd3},
'{3'd3,3'd1,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_15_23[7:0][7:0] = '{'{3'd3,3'd1,3'd0,3'd0,3'd0,3'd1,3'd2,3'd3},
'{3'd3,3'd4,3'd0,3'd0,3'd0,3'd3,3'd3,3'd3},
'{3'd4,3'd0,3'd0,3'd0,3'd4,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3},
'{3'd1,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3},
'{3'd1,3'd0,3'd4,3'd0,3'd1,3'd3,3'd3,3'd3},
'{3'd4,3'd0,3'd0,3'd0,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_15_24[7:0][7:0] = '{'{3'd1,3'd0,3'd0,3'd4,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd0,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_15_25[7:0][7:0] = '{'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd2,3'd3},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd2,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd1,3'd2,3'd3,3'd3,3'd3},
'{3'd0,3'd4,3'd4,3'd0,3'd2,3'd3,3'd2,3'd3},
'{3'd0,3'd4,3'd1,3'd2,3'd3,3'd3,3'd2,3'd2},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_15_26[7:0][7:0] = '{'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd3,3'd3,3'd1,3'd1,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd0,3'd0,3'd4,3'd4,3'd1,3'd1,3'd3},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_15_27[7:0][7:0] = '{'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd2,3'd0,3'd1},
'{3'd0,3'd0,3'd4,3'd4,3'd1,3'd1,3'd0,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd3},
'{3'd0,3'd4,3'd1,3'd0,3'd0,3'd0,3'd3,3'd3},
'{3'd4,3'd4,3'd3,3'd4,3'd0,3'd0,3'd2,3'd3},
'{3'd1,3'd1,3'd3,3'd3,3'd0,3'd0,3'd4,3'd3},
'{3'd1,3'd1,3'd3,3'd3,3'd1,3'd1,3'd1,3'd3},
'{3'd3,3'd3,3'd3,3'd2,3'd2,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_15_28[7:0][7:0] = '{'{3'd3,3'd1,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd1,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd2,3'd1,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3},
'{3'd2,3'd3,3'd2,3'd3,3'd3,3'd3,3'd2,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd2}};

parameter bit [2:0] SpriteTableG_15_29[7:0][7:0] = '{'{3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd1,3'd1},
'{3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1},
'{3'd1,3'd2,3'd2,3'd3,3'd3,3'd3,3'd2,3'd2},
'{3'd2,3'd1,3'd2,3'd3,3'd3,3'd3,3'd2,3'd2},
'{3'd2,3'd4,3'd1,3'd3,3'd3,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0},
'{3'd2,3'd0,3'd0,3'd4,3'd1,3'd4,3'd0,3'd0},
'{3'd3,3'd1,3'd0,3'd3,3'd3,3'd3,3'd0,3'd1}};

parameter bit [2:0] SpriteTableG_15_30[7:0][7:0] = '{'{3'd3,3'd1,3'd0,3'd3,3'd3,3'd3,3'd0,3'd1},
'{3'd3,3'd4,3'd0,3'd1,3'd3,3'd1,3'd0,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd0,3'd0,3'd0,3'd4,3'd0,3'd0,3'd0},
'{3'd3,3'd4,3'd0,3'd1,3'd3,3'd1,3'd0,3'd4},
'{3'd3,3'd1,3'd0,3'd3,3'd3,3'd3,3'd0,3'd1},
'{3'd3,3'd4,3'd0,3'd1,3'd3,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_15_31[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd0,3'd0,3'd2,3'd3,3'd1,3'd0,3'd0},
'{3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd0,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_15_32[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd0},
'{3'd3,3'd3,3'd3,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd2,3'd0,3'd4,3'd3,3'd1,3'd0,3'd0},
'{3'd3,3'd4,3'd0,3'd4,3'd3,3'd4,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_15_33[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd1,3'd4,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd1,3'd4,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_15_34[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_15_35[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_16_0[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_16_1[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd4,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd3,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd3,3'd4,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd4}};

parameter bit [2:0] SpriteTableG_16_2[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd3,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd4,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_16_3[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd4,3'd3,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd4,3'd3,3'd1,3'd0,3'd0,3'd4},
'{3'd0,3'd1,3'd3,3'd1,3'd0,3'd0,3'd0,3'd2},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd1,3'd3},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd3},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd3,3'd3},
'{3'd1,3'd1,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd1,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_16_4[7:0][7:0] = '{'{3'd1,3'd1,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3},
'{3'd1,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3},
'{3'd1,3'd1,3'd0,3'd0,3'd2,3'd3,3'd3,3'd3},
'{3'd1,3'd1,3'd0,3'd0,3'd2,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd0,3'd0,3'd2,3'd1,3'd1,3'd3},
'{3'd1,3'd1,3'd0,3'd0,3'd1,3'd1,3'd3,3'd1},
'{3'd1,3'd1,3'd0,3'd0,3'd4,3'd1,3'd3,3'd1}};

parameter bit [2:0] SpriteTableG_16_5[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd3,3'd4},
'{3'd1,3'd1,3'd0,3'd0,3'd4,3'd3,3'd3,3'd4},
'{3'd3,3'd3,3'd0,3'd0,3'd1,3'd3,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1}};

parameter bit [2:0] SpriteTableG_16_6[7:0][7:0] = '{'{3'd3,3'd3,3'd4,3'd0,3'd1,3'd3,3'd1,3'd1},
'{3'd3,3'd3,3'd4,3'd0,3'd1,3'd3,3'd3,3'd4},
'{3'd1,3'd2,3'd2,3'd0,3'd4,3'd3,3'd1,3'd4},
'{3'd0,3'd2,3'd3,3'd0,3'd4,3'd1,3'd1,3'd4},
'{3'd3,3'd3,3'd3,3'd1,3'd4,3'd1,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0},
'{3'd3,3'd3,3'd3,3'd2,3'd1,3'd3,3'd3,3'd1}};

parameter bit [2:0] SpriteTableG_16_7[7:0][7:0] = '{'{3'd2,3'd2,3'd1,3'd2,3'd3,3'd2,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd3,3'd3,3'd3,3'd2,3'd1},
'{3'd0,3'd0,3'd0,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd0,3'd0,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd1}};

parameter bit [2:0] SpriteTableG_16_8[7:0][7:0] = '{'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd0,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd0,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd0,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4}};

parameter bit [2:0] SpriteTableG_16_9[7:0][7:0] = '{'{3'd0,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0},
'{3'd0,3'd0,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd0,3'd0,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd4,3'd0},
'{3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd0,3'd0},
'{3'd0,3'd4,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0},
'{3'd0,3'd4,3'd3,3'd3,3'd3,3'd1,3'd0,3'd4},
'{3'd0,3'd4,3'd3,3'd3,3'd3,3'd4,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_16_10[7:0][7:0] = '{'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd0,3'd0,3'd4},
'{3'd0,3'd1,3'd3,3'd3,3'd1,3'd0,3'd4,3'd1},
'{3'd0,3'd1,3'd3,3'd3,3'd1,3'd0,3'd0,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd4,3'd0,3'd0,3'd1},
'{3'd0,3'd1,3'd3,3'd1,3'd0,3'd0,3'd4,3'd3},
'{3'd0,3'd1,3'd3,3'd1,3'd0,3'd0,3'd1,3'd3},
'{3'd0,3'd1,3'd3,3'd4,3'd0,3'd0,3'd1,3'd3},
'{3'd0,3'd1,3'd3,3'd0,3'd0,3'd0,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_16_11[7:0][7:0] = '{'{3'd0,3'd1,3'd1,3'd0,3'd4,3'd4,3'd3,3'd3},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd1,3'd3,3'd2},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd3,3'd3,3'd2},
'{3'd0,3'd1,3'd4,3'd0,3'd4,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd0,3'd4,3'd1,3'd3,3'd3,3'd3},
'{3'd0,3'd4,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd2}};

parameter bit [2:0] SpriteTableG_16_12[7:0][7:0] = '{'{3'd0,3'd4,3'd0,3'd1,3'd3,3'd3,3'd2,3'd2},
'{3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_16_13[7:0][7:0] = '{'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_16_14[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_16_15[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_16_16[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd1,3'd1},
'{3'd4,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_16_17[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd1,3'd1,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd4,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd1,3'd4,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_16_18[7:0][7:0] = '{'{3'd3,3'd3,3'd1,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd4,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd1,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd1,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_16_19[7:0][7:0] = '{'{3'd1,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_16_20[7:0][7:0] = '{'{3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_16_21[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_16_22[7:0][7:0] = '{'{3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd2,3'd1,3'd1,3'd0,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd2,3'd1,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_16_23[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd2,3'd2,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd2,3'd0,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_16_24[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd2,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_16_25[7:0][7:0] = '{'{3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd2,3'd3},
'{3'd3,3'd3,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd2,3'd3,3'd2,3'd2,3'd3},
'{3'd3,3'd3,3'd3,3'd2,3'd3,3'd2,3'd2,3'd3},
'{3'd3,3'd3,3'd2,3'd2,3'd3,3'd3,3'd2,3'd3},
'{3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd2,3'd2},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1}};

parameter bit [2:0] SpriteTableG_16_26[7:0][7:0] = '{'{3'd3,3'd1,3'd1,3'd1,3'd4,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4},
'{3'd0,3'd4,3'd1,3'd1,3'd1,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_16_27[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd2,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2}};

parameter bit [2:0] SpriteTableG_16_28[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_16_29[7:0][7:0] = '{'{3'd1,3'd1,3'd2,3'd3,3'd2,3'd2,3'd3,3'd3},
'{3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd3,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd2},
'{3'd3,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd2},
'{3'd3,3'd3,3'd2,3'd1,3'd3,3'd3,3'd3,3'd2},
'{3'd0,3'd1,3'd1,3'd1,3'd3,3'd2,3'd2,3'd2},
'{3'd1,3'd1,3'd0,3'd0,3'd2,3'd3,3'd2,3'd2},
'{3'd3,3'd3,3'd1,3'd0,3'd3,3'd3,3'd3,3'd2}};

parameter bit [2:0] SpriteTableG_16_30[7:0][7:0] = '{'{3'd3,3'd3,3'd1,3'd0,3'd3,3'd3,3'd3,3'd4},
'{3'd3,3'd3,3'd4,3'd0,3'd1,3'd3,3'd2,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd0},
'{3'd4,3'd4,3'd0,3'd0,3'd0,3'd4,3'd0,3'd0},
'{3'd3,3'd3,3'd4,3'd0,3'd1,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd1,3'd0,3'd3,3'd3,3'd3,3'd0},
'{3'd3,3'd3,3'd4,3'd0,3'd1,3'd3,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_16_31[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd3,3'd0,3'd0,3'd4,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd1,3'd0,3'd1,3'd3,3'd3,3'd0},
'{3'd1,3'd3,3'd0,3'd0,3'd4,3'd3,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd4,3'd0},
'{3'd3,3'd3,3'd4,3'd0,3'd1,3'd3,3'd1,3'd0}};

parameter bit [2:0] SpriteTableG_16_32[7:0][7:0] = '{'{3'd1,3'd1,3'd0,3'd0,3'd4,3'd3,3'd4,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd2,3'd4},
'{3'd0,3'd0,3'd0,3'd4,3'd2,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd1,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd3,3'd3,3'd2,3'd3}};

parameter bit [2:0] SpriteTableG_16_33[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd3,3'd1,3'd0,3'd0},
'{3'd4,3'd1,3'd0,3'd0,3'd1,3'd4,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_16_34[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_16_35[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_17_0[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_17_1[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_17_2[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd2,3'd2,3'd1,3'd1,3'd0,3'd0,3'd1,3'd1},
'{3'd1,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd4,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1}};

parameter bit [2:0] SpriteTableG_17_3[7:0][7:0] = '{'{3'd0,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd2,3'd2,3'd1,3'd3,3'd2,3'd1,3'd1,3'd1},
'{3'd3,3'd2,3'd2,3'd3,3'd2,3'd1,3'd1,3'd1},
'{3'd3,3'd2,3'd2,3'd3,3'd2,3'd1,3'd1,3'd1},
'{3'd3,3'd2,3'd2,3'd3,3'd0,3'd1,3'd1,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd1,3'd1}};

parameter bit [2:0] SpriteTableG_17_4[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd0,3'd0,3'd0,3'd1},
'{3'd3,3'd3,3'd3,3'd4,3'd0,3'd0,3'd1,3'd2},
'{3'd3,3'd3,3'd3,3'd0,3'd0,3'd0,3'd1,3'd3},
'{3'd3,3'd3,3'd3,3'd4,3'd0,3'd0,3'd4,3'd1},
'{3'd2,3'd3,3'd3,3'd1,3'd0,3'd0,3'd1,3'd1},
'{3'd0,3'd3,3'd3,3'd1,3'd0,3'd0,3'd1,3'd0},
'{3'd0,3'd3,3'd3,3'd4,3'd0,3'd1,3'd3,3'd1},
'{3'd4,3'd3,3'd1,3'd0,3'd0,3'd1,3'd3,3'd1}};

parameter bit [2:0] SpriteTableG_17_5[7:0][7:0] = '{'{3'd1,3'd1,3'd0,3'd0,3'd4,3'd1,3'd0,3'd0},
'{3'd1,3'd4,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0},
'{3'd1,3'd4,3'd0,3'd0,3'd1,3'd0,3'd4,3'd0},
'{3'd1,3'd1,3'd3,3'd1,3'd1,3'd1,3'd3,3'd1},
'{3'd1,3'd3,3'd3,3'd1,3'd0,3'd1,3'd3,3'd1},
'{3'd1,3'd4,3'd1,3'd1,3'd0,3'd0,3'd1,3'd4},
'{3'd4,3'd0,3'd4,3'd4,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd4,3'd1,3'd0,3'd0,3'd0,3'd1,3'd4}};

parameter bit [2:0] SpriteTableG_17_6[7:0][7:0] = '{'{3'd0,3'd3,3'd3,3'd4,3'd0,3'd1,3'd3,3'd3},
'{3'd4,3'd3,3'd3,3'd1,3'd0,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd4,3'd0,3'd1,3'd3,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd4,3'd1,3'd4},
'{3'd4,3'd3,3'd3,3'd1,3'd0,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd0,3'd3,3'd3,3'd3},
'{3'd4,3'd3,3'd3,3'd1,3'd0,3'd1,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_17_7[7:0][7:0] = '{'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd4,3'd0},
'{3'd1,3'd2,3'd1,3'd4,3'd0,3'd4,3'd1,3'd1},
'{3'd2,3'd3,3'd3,3'd1,3'd0,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd1,3'd4,3'd4,3'd1,3'd4,3'd4},
'{3'd4,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd4,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1}};

parameter bit [2:0] SpriteTableG_17_8[7:0][7:0] = '{'{3'd1,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd0,3'd0,3'd1,3'd3,3'd2,3'd2,3'd2},
'{3'd0,3'd0,3'd0,3'd3,3'd3,3'd2,3'd2,3'd2},
'{3'd0,3'd0,3'd4,3'd3,3'd3,3'd2,3'd2,3'd2},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd2,3'd2,3'd2},
'{3'd0,3'd0,3'd1,3'd3,3'd2,3'd2,3'd2,3'd2},
'{3'd0,3'd0,3'd1,3'd3,3'd2,3'd2,3'd2,3'd2},
'{3'd0,3'd4,3'd3,3'd3,3'd2,3'd3,3'd2,3'd2}};

parameter bit [2:0] SpriteTableG_17_9[7:0][7:0] = '{'{3'd0,3'd4,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd0,3'd1,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd0,3'd1,3'd3,3'd2,3'd2,3'd3,3'd2,3'd2},
'{3'd0,3'd3,3'd3,3'd2,3'd2,3'd3,3'd2,3'd2},
'{3'd4,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd1,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd1,3'd3,3'd3,3'd2,3'd3,3'd3,3'd2,3'd3},
'{3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3}};

parameter bit [2:0] SpriteTableG_17_10[7:0][7:0] = '{'{3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd3},
'{3'd3,3'd2,3'd3,3'd3,3'd2,3'd2,3'd2,3'd3},
'{3'd2,3'd2,3'd2,3'd3,3'd2,3'd2,3'd2,3'd3},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2},
'{3'd2,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd1,3'd2}};

parameter bit [2:0] SpriteTableG_17_11[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd3,3'd2,3'd2,3'd3},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd2,3'd3,3'd2,3'd2,3'd3,3'd2,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2}};

parameter bit [2:0] SpriteTableG_17_12[7:0][7:0] = '{'{3'd3,3'd2,3'd3,3'd3,3'd2,3'd3,3'd2,3'd3},
'{3'd2,3'd3,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_17_13[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_17_14[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd1},
'{3'd2,3'd2,3'd2,3'd3,3'd3,3'd4,3'd0,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd3,3'd3,3'd1,3'd4,3'd0,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd4,3'd0,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd0,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd0,3'd4,3'd0,3'd1}};

parameter bit [2:0] SpriteTableG_17_15[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd4,3'd0,3'd1},
'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd1},
'{3'd3,3'd3,3'd3,3'd4,3'd0,3'd0,3'd0,3'd3},
'{3'd3,3'd3,3'd3,3'd4,3'd0,3'd0,3'd0,3'd3},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd3},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd3},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd4,3'd3},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd4,3'd3}};

parameter bit [2:0] SpriteTableG_17_16[7:0][7:0] = '{'{3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd4,3'd3},
'{3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3},
'{3'd3,3'd1,3'd4,3'd0,3'd0,3'd0,3'd1,3'd3},
'{3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3},
'{3'd0,3'd0,3'd0,3'd4,3'd0,3'd0,3'd4,3'd1},
'{3'd0,3'd0,3'd4,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd4,3'd4,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_17_17[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd4,3'd4,3'd0,3'd1,3'd1,3'd1,3'd3},
'{3'd3,3'd3,3'd3,3'd0,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_17_18[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_17_19[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_17_20[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_17_21[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_17_22[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd1}};

parameter bit [2:0] SpriteTableG_17_23[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd4,3'd0,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd0,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd0,3'd0,3'd4,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd0,3'd0,3'd1,3'd3},
'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd1,3'd3},
'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd1,3'd1},
'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_17_24[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd4,3'd4,3'd1,3'd0,3'd4},
'{3'd3,3'd3,3'd3,3'd0,3'd0,3'd4,3'd4,3'd1},
'{3'd3,3'd3,3'd1,3'd1,3'd1,3'd3,3'd3,3'd3},
'{3'd3,3'd1,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd2,3'd3,3'd3,3'd2,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3},
'{3'd2,3'd2,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_17_25[7:0][7:0] = '{'{3'd3,3'd3,3'd2,3'd3,3'd3,3'd2,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3},
'{3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd0,3'd0,3'd4,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_17_26[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_17_27[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd3,3'd3,3'd2,3'd2,3'd3,3'd3,3'd3},
'{3'd1,3'd2,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_17_28[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd2,3'd1,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd2,3'd1,3'd1,3'd1,3'd2,3'd1},
'{3'd3,3'd3,3'd3,3'd2,3'd1,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_17_29[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd2,3'd3,3'd3,3'd2,3'd1,3'd2,3'd3,3'd2},
'{3'd2,3'd3,3'd3,3'd3,3'd1,3'd3,3'd3,3'd3},
'{3'd2,3'd3,3'd3,3'd1,3'd0,3'd3,3'd3,3'd3},
'{3'd2,3'd3,3'd3,3'd4,3'd0,3'd2,3'd3,3'd2},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd2,3'd1},
'{3'd4,3'd3,3'd3,3'd1,3'd0,3'd1,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_17_30[7:0][7:0] = '{'{3'd1,3'd3,3'd3,3'd1,3'd0,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd4,3'd0,3'd1,3'd3,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd0,3'd3,3'd3,3'd4,3'd0,3'd4,3'd3,3'd2},
'{3'd4,3'd3,3'd3,3'd1,3'd0,3'd1,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd4,3'd0,3'd4,3'd3,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_17_31[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd4,3'd1,3'd1},
'{3'd0,3'd3,3'd3,3'd1,3'd0,3'd1,3'd3,3'd1},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd4,3'd1,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd4,3'd4,3'd0,3'd0,3'd0,3'd4,3'd0},
'{3'd0,3'd3,3'd3,3'd0,3'd0,3'd4,3'd3,3'd1}};

parameter bit [2:0] SpriteTableG_17_32[7:0][7:0] = '{'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd4},
'{3'd1,3'd4,3'd1,3'd0,3'd0,3'd0,3'd1,3'd0},
'{3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_17_33[7:0][7:0] = '{'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_17_34[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd2,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_17_35[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_18_0[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_18_1[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_18_2[7:0][7:0] = '{'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd2,3'd1,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd2,3'd3,3'd3,3'd1,3'd0},
'{3'd1,3'd1,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd1,3'd1,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd1,3'd1,3'd3,3'd3,3'd3,3'd3,3'd2}};

parameter bit [2:0] SpriteTableG_18_3[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd3,3'd2,3'd1,3'd3,3'd3},
'{3'd1,3'd1,3'd2,3'd3,3'd1,3'd1,3'd2,3'd3},
'{3'd1,3'd1,3'd3,3'd2,3'd2,3'd3,3'd3,3'd2},
'{3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd2,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2}};

parameter bit [2:0] SpriteTableG_18_4[7:0][7:0] = '{'{3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2},
'{3'd1,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1},
'{3'd4,3'd0,3'd4,3'd1,3'd0,3'd0,3'd0,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd4,3'd0,3'd0,3'd0,3'd4},
'{3'd0,3'd0,3'd1,3'd3,3'd0,3'd0,3'd4,3'd3},
'{3'd0,3'd0,3'd1,3'd3,3'd0,3'd0,3'd4,3'd3}};

parameter bit [2:0] SpriteTableG_18_5[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd4,3'd1,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd4,3'd3,3'd3,3'd1,3'd0,3'd1,3'd3},
'{3'd0,3'd4,3'd3,3'd3,3'd1,3'd0,3'd1,3'd3},
'{3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd4,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1}};

parameter bit [2:0] SpriteTableG_18_6[7:0][7:0] = '{'{3'd0,3'd4,3'd3,3'd3,3'd1,3'd0,3'd1,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd1,3'd0,3'd3,3'd3},
'{3'd0,3'd0,3'd3,3'd3,3'd1,3'd0,3'd1,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd4,3'd2},
'{3'd0,3'd1,3'd3,3'd3,3'd1,3'd0,3'd3,3'd3},
'{3'd4,3'd1,3'd3,3'd3,3'd3,3'd4,3'd3,3'd3},
'{3'd0,3'd4,3'd3,3'd3,3'd1,3'd0,3'd1,3'd3}};

parameter bit [2:0] SpriteTableG_18_7[7:0][7:0] = '{'{3'd0,3'd0,3'd4,3'd4,3'd0,3'd0,3'd1,3'd0},
'{3'd0,3'd0,3'd1,3'd1,3'd4,3'd1,3'd0,3'd0},
'{3'd4,3'd1,3'd3,3'd3,3'd2,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd3,3'd2,3'd1,3'd1,3'd1,3'd1},
'{3'd4,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd1},
'{3'd1,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_18_8[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd3,3'd2,3'd2,3'd3,3'd2,3'd2,3'd3,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd3,3'd2,3'd2,3'd3,3'd2,3'd2,3'd3,3'd2}};

parameter bit [2:0] SpriteTableG_18_9[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd3,3'd2,3'd2,3'd3,3'd2,3'd2,3'd3,3'd2},
'{3'd3,3'd2,3'd2,3'd3,3'd2,3'd2,3'd3,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd3,3'd2,3'd3,3'd3,3'd2,3'd3,3'd3,3'd2},
'{3'd3,3'd2,3'd2,3'd3,3'd2,3'd2,3'd3,3'd2}};

parameter bit [2:0] SpriteTableG_18_10[7:0][7:0] = '{'{3'd2,3'd3,3'd2,3'd2,3'd3,3'd2,3'd2,3'd2},
'{3'd3,3'd2,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3},
'{3'd3,3'd2,3'd3,3'd3,3'd2,3'd3,3'd3,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd2,3'd3},
'{3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_18_11[7:0][7:0] = '{'{3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_18_12[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_18_13[7:0][7:0] = '{'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_18_14[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd1,3'd1,3'd2,3'd2,3'd2,3'd3,3'd3},
'{3'd4,3'd0,3'd4,3'd1,3'd1,3'd1,3'd1,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_18_15[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_18_16[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd4,3'd4,3'd4,3'd0},
'{3'd0,3'd0,3'd0,3'd4,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_18_17[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd4,3'd4,3'd4,3'd1,3'd1,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2}};

parameter bit [2:0] SpriteTableG_18_18[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd1},
'{3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_18_19[7:0][7:0] = '{'{3'd3,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd0,3'd0,3'd4,3'd1,3'd1,3'd1,3'd1},
'{3'd3,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd0,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd0,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_18_20[7:0][7:0] = '{'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd4,3'd1,3'd0,3'd0,3'd4,3'd0},
'{3'd1,3'd0,3'd4,3'd1,3'd4,3'd1,3'd1,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_18_21[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_18_22[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd4,3'd4,3'd4,3'd4,3'd4,3'd4,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1}};

parameter bit [2:0] SpriteTableG_18_23[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd4,3'd4,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_18_24[7:0][7:0] = '{'{3'd1,3'd0,3'd4,3'd1,3'd1,3'd1,3'd3,3'd0},
'{3'd1,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd4},
'{3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1}};

parameter bit [2:0] SpriteTableG_18_25[7:0][7:0] = '{'{3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd1,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd1,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd3},
'{3'd3,3'd1,3'd1,3'd1,3'd1,3'd4,3'd1,3'd3},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd4,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_18_26[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd3},
'{3'd1,3'd3,3'd1,3'd0,3'd0,3'd4,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd0,3'd0,3'd0,3'd4,3'd0},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd1,3'd2},
'{3'd3,3'd3,3'd1,3'd1,3'd3,3'd0,3'd0,3'd3},
'{3'd1,3'd1,3'd3,3'd3,3'd3,3'd2,3'd2,3'd3}};

parameter bit [2:0] SpriteTableG_18_27[7:0][7:0] = '{'{3'd0,3'd1,3'd3,3'd3,3'd2,3'd1,3'd2,3'd3},
'{3'd1,3'd1,3'd3,3'd3,3'd2,3'd1,3'd2,3'd3},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd1,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3},
'{3'd1,3'd1,3'd3,3'd3,3'd2,3'd1,3'd2,3'd3},
'{3'd1,3'd1,3'd2,3'd2,3'd1,3'd1,3'd1,3'd2},
'{3'd2,3'd2,3'd3,3'd3,3'd3,3'd1,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_18_28[7:0][7:0] = '{'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3},
'{3'd2,3'd2,3'd3,3'd3,3'd3,3'd1,3'd3,3'd3},
'{3'd2,3'd2,3'd3,3'd3,3'd2,3'd1,3'd2,3'd3},
'{3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd2,3'd2,3'd3,3'd3,3'd2,3'd1,3'd2,3'd3},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd1,3'd3,3'd3},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd1,3'd3,3'd3},
'{3'd1,3'd1,3'd3,3'd3,3'd2,3'd1,3'd2,3'd3}};

parameter bit [2:0] SpriteTableG_18_29[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd2,3'd3,3'd1,3'd1,3'd1,3'd3},
'{3'd1,3'd2,3'd3,3'd3,3'd3,3'd0,3'd1,3'd3},
'{3'd1,3'd2,3'd3,3'd3,3'd1,3'd0,3'd3,3'd3},
'{3'd1,3'd1,3'd3,3'd3,3'd1,3'd0,3'd4,3'd3},
'{3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd2,3'd2,3'd0,3'd0,3'd0,3'd4},
'{3'd1,3'd1,3'd3,3'd3,3'd1,3'd0,3'd1,3'd3}};

parameter bit [2:0] SpriteTableG_18_30[7:0][7:0] = '{'{3'd2,3'd2,3'd3,3'd3,3'd1,3'd0,3'd1,3'd3},
'{3'd1,3'd1,3'd2,3'd1,3'd4,3'd0,3'd4,3'd1},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd3,3'd4,3'd0,3'd4,3'd1},
'{3'd0,3'd0,3'd3,3'd3,3'd1,3'd0,3'd1,3'd3},
'{3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_18_31[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd3,3'd3,3'd4,3'd0,3'd4,3'd3},
'{3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd3,3'd0,3'd0,3'd0,3'd1}};

parameter bit [2:0] SpriteTableG_18_32[7:0][7:0] = '{'{3'd0,3'd0,3'd4,3'd1,3'd0,3'd0,3'd0,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_18_33[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd2,3'd4,3'd1,3'd1,3'd2,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_18_34[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0},
'{3'd3,3'd3,3'd2,3'd0,3'd1,3'd1,3'd2,3'd1},
'{3'd3,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_18_35[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_19_0[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_19_1[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_19_2[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd2,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd4,3'd2,3'd3,3'd1,3'd0,3'd0},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd4,3'd0,3'd0},
'{3'd2,3'd3,3'd3,3'd2,3'd2,3'd4,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_19_3[7:0][7:0] = '{'{3'd3,3'd3,3'd2,3'd2,3'd3,3'd4,3'd0,3'd0},
'{3'd3,3'd3,3'd2,3'd2,3'd3,3'd3,3'd4,3'd0},
'{3'd2,3'd3,3'd3,3'd2,3'd2,3'd3,3'd3,3'd4},
'{3'd2,3'd3,3'd3,3'd3,3'd2,3'd2,3'd3,3'd3},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1},
'{3'd2,3'd3,3'd3,3'd3,3'd1,3'd4,3'd0,3'd0},
'{3'd2,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_19_4[7:0][7:0] = '{'{3'd2,3'd3,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd2,3'd4,3'd1,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd2,3'd1,3'd2,3'd0,3'd0,3'd0},
'{3'd2,3'd3,3'd2,3'd2,3'd1,3'd1,3'd1,3'd4},
'{3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1},
'{3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1},
'{3'd1,3'd1,3'd2,3'd3,3'd3,3'd2,3'd1,3'd2},
'{3'd1,3'd1,3'd2,3'd3,3'd3,3'd2,3'd1,3'd2}};

parameter bit [2:0] SpriteTableG_19_5[7:0][7:0] = '{'{3'd0,3'd0,3'd2,3'd2,3'd2,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd1,3'd2,3'd1,3'd2,3'd1,3'd1},
'{3'd4,3'd0,3'd1,3'd2,3'd3,3'd2,3'd1,3'd1},
'{3'd3,3'd0,3'd2,3'd3,3'd3,3'd2,3'd1,3'd3},
'{3'd3,3'd0,3'd1,3'd3,3'd3,3'd3,3'd1,3'd3},
'{3'd1,3'd0,3'd1,3'd2,3'd3,3'd2,3'd1,3'd2},
'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd4,3'd0,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1}};

parameter bit [2:0] SpriteTableG_19_6[7:0][7:0] = '{'{3'd3,3'd1,3'd2,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd3,3'd2,3'd2,3'd3,3'd3,3'd2,3'd0,3'd1},
'{3'd3,3'd2,3'd2,3'd3,3'd2,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd1,3'd0},
'{3'd3,3'd2,3'd1,3'd0,3'd0,3'd0,3'd1,3'd0},
'{3'd3,3'd2,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0},
'{3'd3,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1}};

parameter bit [2:0] SpriteTableG_19_7[7:0][7:0] = '{'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd0},
'{3'd1,3'd1,3'd1,3'd3,3'd3,3'd3,3'd3,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0}};

parameter bit [2:0] SpriteTableG_19_8[7:0][7:0] = '{'{3'd2,3'd3,3'd2,3'd2,3'd2,3'd3,3'd3,3'd0},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd0},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd1,3'd0},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd1,3'd0},
'{3'd2,3'd3,3'd2,3'd2,3'd3,3'd3,3'd1,3'd0},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd1,3'd0},
'{3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd4,3'd0},
'{3'd2,3'd3,3'd2,3'd2,3'd3,3'd3,3'd4,3'd0}};

parameter bit [2:0] SpriteTableG_19_9[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd0,3'd0},
'{3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd0,3'd0},
'{3'd2,3'd3,3'd2,3'd2,3'd3,3'd1,3'd0,3'd0},
'{3'd2,3'd3,3'd2,3'd2,3'd3,3'd1,3'd0,3'd0},
'{3'd2,3'd2,3'd2,3'd2,3'd3,3'd1,3'd0,3'd0},
'{3'd2,3'd2,3'd2,3'd2,3'd3,3'd1,3'd0,3'd0},
'{3'd3,3'd3,3'd2,3'd3,3'd3,3'd4,3'd0,3'd4},
'{3'd2,3'd3,3'd2,3'd3,3'd3,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_19_10[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd3,3'd3,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd2,3'd3,3'd3,3'd0,3'd0,3'd1},
'{3'd3,3'd3,3'd2,3'd3,3'd1,3'd0,3'd0,3'd1},
'{3'd2,3'd3,3'd2,3'd3,3'd1,3'd0,3'd0,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd4,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd1,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd1,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd0,3'd0,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_19_11[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd1,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd4,3'd1,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd1,3'd1,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd4,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd1,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_19_12[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd1,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd3}};

parameter bit [2:0] SpriteTableG_19_13[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_19_14[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_19_15[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0},
'{3'd3,3'd1,3'd1,3'd3,3'd3,3'd4,3'd0,3'd0},
'{3'd3,3'd3,3'd1,3'd1,3'd3,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd1,3'd4,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd1,3'd4,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_19_16[7:0][7:0] = '{'{3'd1,3'd3,3'd3,3'd0,3'd0,3'd4,3'd4,3'd0},
'{3'd0,3'd3,3'd1,3'd0,3'd0,3'd1,3'd4,3'd0},
'{3'd4,3'd3,3'd1,3'd0,3'd0,3'd1,3'd4,3'd0},
'{3'd1,3'd3,3'd4,3'd0,3'd0,3'd3,3'd4,3'd0},
'{3'd3,3'd1,3'd0,3'd0,3'd1,3'd3,3'd4,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_19_17[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd1},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd3},
'{3'd2,3'd3,3'd3,3'd2,3'd2,3'd3,3'd2,3'd3},
'{3'd3,3'd3,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd3,3'd3,3'd2,3'd2,3'd3,3'd3,3'd1},
'{3'd2,3'd3,3'd3,3'd3,3'd2,3'd2,3'd3,3'd1}};

parameter bit [2:0] SpriteTableG_19_18[7:0][7:0] = '{'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0},
'{3'd2,3'd3,3'd2,3'd2,3'd2,3'd3,3'd1,3'd4},
'{3'd2,3'd3,3'd3,3'd2,3'd2,3'd3,3'd4,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd1},
'{3'd4,3'd4,3'd4,3'd4,3'd4,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1}};

parameter bit [2:0] SpriteTableG_19_19[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd4,3'd0,3'd0,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd0,3'd3},
'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd4,3'd3},
'{3'd3,3'd4,3'd4,3'd4,3'd0,3'd0,3'd1,3'd3},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3},
'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_19_20[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd0,3'd4,3'd0,3'd0,3'd4,3'd1,3'd3,3'd3},
'{3'd1,3'd1,3'd4,3'd0,3'd4,3'd1,3'd3,3'd3},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd4,3'd0,3'd4,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_19_21[7:0][7:0] = '{'{3'd3,3'd3,3'd4,3'd0,3'd1,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd0,3'd0,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd0,3'd0,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd1,3'd0,3'd0,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd1,3'd0,3'd4,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd1,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_19_22[7:0][7:0] = '{'{3'd3,3'd4,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd4,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_19_23[7:0][7:0] = '{'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_19_24[7:0][7:0] = '{'{3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_19_25[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd1}};

parameter bit [2:0] SpriteTableG_19_26[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd1,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd0,3'd0,3'd0,3'd4,3'd1,3'd1,3'd3,3'd3},
'{3'd4,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd0}};

parameter bit [2:0] SpriteTableG_19_27[7:0][7:0] = '{'{3'd3,3'd2,3'd1,3'd2,3'd3,3'd3,3'd2,3'd0},
'{3'd2,3'd0,3'd0,3'd0,3'd1,3'd3,3'd2,3'd0},
'{3'd3,3'd2,3'd1,3'd0,3'd0,3'd1,3'd1,3'd0},
'{3'd3,3'd1,3'd2,3'd2,3'd0,3'd1,3'd0,3'd0},
'{3'd3,3'd1,3'd1,3'd3,3'd2,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd1,3'd3,3'd1,3'd1,3'd0},
'{3'd4,3'd0,3'd0,3'd4,3'd4,3'd0,3'd1,3'd1},
'{3'd3,3'd4,3'd4,3'd3,3'd3,3'd1,3'd0,3'd2}};

parameter bit [2:0] SpriteTableG_19_28[7:0][7:0] = '{'{3'd3,3'd1,3'd1,3'd3,3'd3,3'd3,3'd4,3'd3},
'{3'd3,3'd2,3'd1,3'd3,3'd3,3'd3,3'd0,3'd3},
'{3'd2,3'd1,3'd1,3'd2,3'd3,3'd4,3'd0,3'd4},
'{3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd1,3'd1,3'd3,3'd3,3'd1,3'd0,3'd4},
'{3'd3,3'd2,3'd2,3'd3,3'd3,3'd3,3'd0,3'd3},
'{3'd3,3'd2,3'd2,3'd3,3'd3,3'd3,3'd1,3'd3},
'{3'd3,3'd1,3'd1,3'd2,3'd3,3'd4,3'd0,3'd4}};

parameter bit [2:0] SpriteTableG_19_29[7:0][7:0] = '{'{3'd1,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd1,3'd4,3'd1,3'd1,3'd4,3'd0,3'd0},
'{3'd3,3'd4,3'd4,3'd3,3'd3,3'd1,3'd0,3'd1},
'{3'd3,3'd4,3'd4,3'd3,3'd3,3'd1,3'd0,3'd1},
'{3'd1,3'd0,3'd0,3'd1,3'd1,3'd4,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd0,3'd0,3'd1},
'{3'd3,3'd4,3'd0,3'd1,3'd3,3'd1,3'd1,3'd1}};

parameter bit [2:0] SpriteTableG_19_30[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd2},
'{3'd4,3'd1,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2},
'{3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd0,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_19_31[7:0][7:0] = '{'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_19_32[7:0][7:0] = '{'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_19_33[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_19_34[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_19_35[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_20_0[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_20_1[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd1,3'd1}};

parameter bit [2:0] SpriteTableG_20_2[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_20_3[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1}};

parameter bit [2:0] SpriteTableG_20_4[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1},
'{3'd3,3'd1,3'd0,3'd0,3'd2,3'd2,3'd1,3'd1},
'{3'd1,3'd4,3'd0,3'd1,3'd2,3'd2,3'd1,3'd1},
'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd2,3'd2,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1},
'{3'd3,3'd3,3'd2,3'd2,3'd3,3'd3,3'd2,3'd1},
'{3'd3,3'd3,3'd2,3'd2,3'd3,3'd3,3'd2,3'd0}};

parameter bit [2:0] SpriteTableG_20_5[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd0,3'd0},
'{3'd1,3'd1,3'd2,3'd2,3'd2,3'd0,3'd1,3'd0},
'{3'd2,3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd2,3'd1,3'd0,3'd1,3'd0,3'd1},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd3,3'd2,3'd0,3'd1,3'd0,3'd1,3'd1,3'd1},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_20_6[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd0,3'd0,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd0,3'd3,3'd3,3'd3,3'd3,3'd4},
'{3'd1,3'd0,3'd2,3'd3,3'd3,3'd3,3'd4,3'd0},
'{3'd0,3'd2,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_20_7[7:0][7:0] = '{'{3'd2,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd4,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd3,3'd3,3'd4,3'd0,3'd0,3'd4},
'{3'd0,3'd4,3'd3,3'd1,3'd0,3'd0,3'd4,3'd3},
'{3'd0,3'd4,3'd3,3'd1,3'd0,3'd0,3'd1,3'd3}};

parameter bit [2:0] SpriteTableG_20_8[7:0][7:0] = '{'{3'd0,3'd1,3'd3,3'd0,3'd0,3'd4,3'd3,3'd3},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd1,3'd3,3'd2},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd3,3'd3,3'd2},
'{3'd0,3'd1,3'd0,3'd0,3'd4,3'd3,3'd3,3'd2},
'{3'd0,3'd4,3'd0,3'd0,3'd1,3'd3,3'd2,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd3,3'd3,3'd2,3'd2},
'{3'd0,3'd0,3'd0,3'd4,3'd3,3'd3,3'd2,3'd2},
'{3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd2,3'd2}};

parameter bit [2:0] SpriteTableG_20_9[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd3,3'd3,3'd2,3'd2,3'd2},
'{3'd0,3'd0,3'd4,3'd3,3'd2,3'd2,3'd2,3'd2},
'{3'd0,3'd0,3'd1,3'd3,3'd2,3'd3,3'd2,3'd2},
'{3'd0,3'd0,3'd3,3'd3,3'd2,3'd3,3'd2,3'd2},
'{3'd0,3'd1,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd0,3'd1,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd0,3'd3,3'd3,3'd2,3'd2,3'd3,3'd2,3'd2},
'{3'd1,3'd3,3'd3,3'd2,3'd2,3'd3,3'd2,3'd2}};

parameter bit [2:0] SpriteTableG_20_10[7:0][7:0] = '{'{3'd1,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3,3'd2},
'{3'd3,3'd2,3'd2,3'd3,3'd3,3'd2,3'd3,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_20_11[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_20_12[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd2,3'd3},
'{3'd3,3'd3,3'd3,3'd4,3'd0,3'd0,3'd1,3'd3},
'{3'd3,3'd3,3'd3,3'd4,3'd0,3'd0,3'd1,3'd3},
'{3'd3,3'd3,3'd3,3'd1,3'd1,3'd2,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd1,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_20_13[7:0][7:0] = '{'{3'd3,3'd3,3'd1,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd1,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd1,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd4,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_20_14[7:0][7:0] = '{'{3'd4,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_20_15[7:0][7:0] = '{'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_20_16[7:0][7:0] = '{'{3'd0,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2},
'{3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd3,3'd3,3'd1,3'd1,3'd1,3'd4,3'd0},
'{3'd0,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd4}};

parameter bit [2:0] SpriteTableG_20_17[7:0][7:0] = '{'{3'd1,3'd0,3'd0,3'd0,3'd4,3'd4,3'd0,3'd0},
'{3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd4,3'd0,3'd0,3'd4,3'd1,3'd3,3'd3,3'd3},
'{3'd4,3'd1,3'd3,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd2,3'd2,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_20_18[7:0][7:0] = '{'{3'd1,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd2},
'{3'd1,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd2},
'{3'd3,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_20_19[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_20_20[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_20_21[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_20_22[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_20_23[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1}};

parameter bit [2:0] SpriteTableG_20_24[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0}};

parameter bit [2:0] SpriteTableG_20_25[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd4,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd4,3'd0,3'd4},
'{3'd4,3'd0,3'd4,3'd0,3'd0,3'd0,3'd0,3'd1}};

parameter bit [2:0] SpriteTableG_20_26[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd1,3'd3},
'{3'd0,3'd0,3'd4,3'd1,3'd3,3'd3,3'd1,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd1},
'{3'd4,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0},
'{3'd1,3'd0,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0},
'{3'd3,3'd1,3'd4,3'd2,3'd3,3'd3,3'd0,3'd0},
'{3'd2,3'd1,3'd0,3'd0,3'd3,3'd3,3'd4,3'd0},
'{3'd0,3'd0,3'd1,3'd0,3'd1,3'd3,3'd1,3'd0}};

parameter bit [2:0] SpriteTableG_20_27[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd1,3'd0,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd0,3'd0,3'd1,3'd1,3'd0,3'd1},
'{3'd0,3'd0,3'd1,3'd0,3'd3,3'd3,3'd3,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd3,3'd3,3'd3,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd2,3'd1,3'd4,3'd1},
'{3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd1,3'd0,3'd1,3'd0,3'd3,3'd3,3'd2,3'd1}};

parameter bit [2:0] SpriteTableG_20_28[7:0][7:0] = '{'{3'd3,3'd1,3'd0,3'd1,3'd3,3'd3,3'd3,3'd0},
'{3'd3,3'd3,3'd1,3'd0,3'd3,3'd3,3'd1,3'd0},
'{3'd1,3'd1,3'd4,3'd1,3'd2,3'd1,3'd4,3'd0},
'{3'd0,3'd4,3'd4,3'd0,3'd1,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd4,3'd0,3'd1,3'd3,3'd4,3'd2},
'{3'd3,3'd3,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd1,3'd4,3'd0,3'd1,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_20_29[7:0][7:0] = '{'{3'd0,3'd1,3'd4,3'd0,3'd1,3'd2,3'd1,3'd2},
'{3'd1,3'd1,3'd4,3'd0,3'd1,3'd1,3'd0,3'd1},
'{3'd3,3'd3,3'd4,3'd0,3'd3,3'd3,3'd1,3'd1},
'{3'd3,3'd3,3'd4,3'd0,3'd3,3'd3,3'd1,3'd4},
'{3'd2,3'd3,3'd4,3'd0,3'd2,3'd3,3'd4,3'd4},
'{3'd1,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd0},
'{3'd1,3'd3,3'd2,3'd2,3'd2,3'd1,3'd1,3'd0},
'{3'd3,3'd3,3'd2,3'd1,3'd1,3'd3,3'd1,3'd0}};

parameter bit [2:0] SpriteTableG_20_30[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd1,3'd1,3'd3,3'd3,3'd0},
'{3'd2,3'd3,3'd2,3'd2,3'd2,3'd1,3'd3,3'd4},
'{3'd2,3'd3,3'd3,3'd2,3'd3,3'd4,3'd3,3'd4},
'{3'd2,3'd3,3'd3,3'd2,3'd1,3'd1,3'd1,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd1,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_20_31[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd3},
'{3'd3,3'd3,3'd3,3'd2,3'd1,3'd3,3'd0,3'd3},
'{3'd3,3'd3,3'd3,3'd0,3'd4,3'd3,3'd0,3'd3},
'{3'd3,3'd3,3'd2,3'd0,3'd0,3'd3,3'd0,3'd1},
'{3'd3,3'd3,3'd2,3'd0,3'd0,3'd3,3'd4,3'd1},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd4,3'd0,3'd0,3'd3,3'd1,3'd0},
'{3'd1,3'd3,3'd0,3'd0,3'd0,3'd3,3'd1,3'd0}};

parameter bit [2:0] SpriteTableG_20_32[7:0][7:0] = '{'{3'd1,3'd3,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0},
'{3'd1,3'd3,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0},
'{3'd1,3'd3,3'd0,3'd0,3'd0,3'd1,3'd3,3'd0},
'{3'd1,3'd3,3'd0,3'd0,3'd0,3'd1,3'd3,3'd0},
'{3'd1,3'd3,3'd0,3'd0,3'd0,3'd1,3'd3,3'd0},
'{3'd1,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1}};

parameter bit [2:0] SpriteTableG_20_33[7:0][7:0] = '{'{3'd3,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3},
'{3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd2,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd3},
'{3'd0,3'd0,3'd0,3'd4,3'd4,3'd0,3'd0,3'd4},
'{3'd0,3'd0,3'd0,3'd4,3'd0,3'd0,3'd4,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_20_34[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd3,3'd2}};

parameter bit [2:0] SpriteTableG_20_35[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd4,3'd2,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd2,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd2,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_21_0[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_21_1[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_21_2[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_21_3[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1}};

parameter bit [2:0] SpriteTableG_21_4[7:0][7:0] = '{'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0},
'{3'd1,3'd2,3'd1,3'd0,3'd1,3'd1,3'd1,3'd0},
'{3'd1,3'd2,3'd4,3'd1,3'd0,3'd0,3'd1,3'd0},
'{3'd1,3'd1,3'd1,3'd0,3'd1,3'd0,3'd1,3'd0},
'{3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1,3'd2},
'{3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd2,3'd3},
'{3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd2,3'd3},
'{3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd2,3'd3}};

parameter bit [2:0] SpriteTableG_21_5[7:0][7:0] = '{'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd2,3'd3},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd3},
'{3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd2,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd2,3'd1,3'd0,3'd2,3'd2},
'{3'd0,3'd0,3'd3,3'd3,3'd0,3'd0,3'd1,3'd1},
'{3'd0,3'd3,3'd3,3'd3,3'd0,3'd0,3'd1,3'd3}};

parameter bit [2:0] SpriteTableG_21_6[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd0,3'd0,3'd2,3'd3},
'{3'd3,3'd3,3'd3,3'd2,3'd0,3'd0,3'd0,3'd3},
'{3'd3,3'd3,3'd3,3'd2,3'd0,3'd0,3'd0,3'd3},
'{3'd3,3'd3,3'd3,3'd2,3'd0,3'd0,3'd0,3'd2},
'{3'd1,3'd3,3'd3,3'd2,3'd0,3'd1,3'd0,3'd1},
'{3'd1,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd3,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_21_7[7:0][7:0] = '{'{3'd1,3'd3,3'd3,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd1,3'd3,3'd3,3'd1,3'd1,3'd1,3'd1,3'd0},
'{3'd4,3'd4,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableG_21_8[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd3,3'd2,3'd2,3'd3,3'd2,3'd2,3'd3,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd3,3'd2,3'd2,3'd3,3'd2,3'd2,3'd3,3'd2}};

parameter bit [2:0] SpriteTableG_21_9[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd3,3'd2,3'd2,3'd3,3'd2,3'd2,3'd3,3'd2},
'{3'd3,3'd2,3'd2,3'd3,3'd2,3'd2,3'd3,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd3,3'd2,3'd2,3'd3,3'd2,3'd2,3'd3,3'd2},
'{3'd3,3'd2,3'd2,3'd3,3'd2,3'd2,3'd3,3'd3},
'{3'd3,3'd2,3'd2,3'd3,3'd2,3'd2,3'd3,3'd2}};

parameter bit [2:0] SpriteTableG_21_10[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd2,3'd3,3'd3,3'd3,3'd2,3'd3},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_21_11[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_21_12[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_21_13[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_21_14[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd3,3'd3},
'{3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_21_15[7:0][7:0] = '{'{3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_21_16[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd3,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd0},
'{3'd4,3'd4,3'd4,3'd1,3'd1,3'd1,3'd4,3'd0},
'{3'd4,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_21_17[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd1,3'd1},
'{3'd1,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_21_18[7:0][7:0] = '{'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd3},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd3},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3},
'{3'd2,3'd2,3'd3,3'd3,3'd2,3'd2,3'd3,3'd3},
'{3'd3,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_21_19[7:0][7:0] = '{'{3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd1,3'd1},
'{3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd0,3'd0},
'{3'd2,3'd2,3'd3,3'd3,3'd3,3'd1,3'd4,3'd4},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd0,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd0,3'd4}};

parameter bit [2:0] SpriteTableG_21_20[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd0,3'd0,3'd1,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd1,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_21_21[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd4,3'd0,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_21_22[7:0][7:0] = '{'{3'd3,3'd3,3'd2,3'd1,3'd2,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_21_23[7:0][7:0] = '{'{3'd1,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_21_24[7:0][7:0] = '{'{3'd4,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd4,3'd1,3'd3,3'd3,3'd3},
'{3'd0,3'd4,3'd0,3'd4,3'd1,3'd3,3'd3,3'd2},
'{3'd0,3'd1,3'd4,3'd0,3'd4,3'd3,3'd2,3'd0},
'{3'd0,3'd1,3'd0,3'd0,3'd0,3'd3,3'd3,3'd3},
'{3'd4,3'd3,3'd1,3'd0,3'd0,3'd1,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_21_25[7:0][7:0] = '{'{3'd4,3'd3,3'd3,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd4,3'd0,3'd0,3'd3,3'd2},
'{3'd1,3'd3,3'd3,3'd1,3'd0,3'd4,3'd1,3'd0},
'{3'd1,3'd3,3'd3,3'd1,3'd0,3'd4,3'd4,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd0,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd1,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd1}};

parameter bit [2:0] SpriteTableG_21_26[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd0,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0},
'{3'd3,3'd3,3'd1,3'd4,3'd0,3'd4,3'd0,3'd0},
'{3'd1,3'd3,3'd1,3'd0,3'd0,3'd1,3'd1,3'd4},
'{3'd1,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_21_27[7:0][7:0] = '{'{3'd1,3'd2,3'd3,3'd2,3'd2,3'd2,3'd3,3'd3},
'{3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3},
'{3'd2,3'd3,3'd3,3'd2,3'd2,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd2,3'd2,3'd3,3'd3,3'd3},
'{3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3},
'{3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd3,3'd3},
'{3'd2,3'd3,3'd3,3'd2,3'd2,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_21_28[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd2,3'd2,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd2,3'd2,3'd3,3'd3,3'd3},
'{3'd4,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_21_29[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd3},
'{3'd1,3'd3,3'd1,3'd0,3'd0,3'd1,3'd3,3'd2},
'{3'd1,3'd3,3'd3,3'd0,3'd0,3'd1,3'd3,3'd4},
'{3'd1,3'd4,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd3,3'd4,3'd0,3'd0,3'd4,3'd1,3'd0}};

parameter bit [2:0] SpriteTableG_21_30[7:0][7:0] = '{'{3'd4,3'd3,3'd1,3'd0,3'd0,3'd4,3'd1,3'd0},
'{3'd0,3'd1,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd4,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd3,3'd1,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd1,3'd1},
'{3'd1,3'd0,3'd1,3'd3,3'd0,3'd0,3'd1,3'd1}};

parameter bit [2:0] SpriteTableG_21_31[7:0][7:0] = '{'{3'd4,3'd0,3'd0,3'd3,3'd4,3'd0,3'd0,3'd1},
'{3'd1,3'd0,3'd0,3'd3,3'd1,3'd0,3'd0,3'd1},
'{3'd1,3'd0,3'd0,3'd1,3'd3,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd1,3'd3,3'd0,3'd0,3'd0},
'{3'd3,3'd0,3'd0,3'd0,3'd3,3'd1,3'd0,3'd0},
'{3'd4,3'd0,3'd0,3'd0,3'd3,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd1,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_21_32[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd4,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_21_33[7:0][7:0] = '{'{3'd2,3'd1,3'd1,3'd2,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd2,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd2,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd4,3'd0,3'd0},
'{3'd2,3'd3,3'd2,3'd1,3'd1,3'd4,3'd0,3'd0},
'{3'd2,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd1,3'd3,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2}};

parameter bit [2:0] SpriteTableG_21_34[7:0][7:0] = '{'{3'd1,3'd3,3'd3,3'd1,3'd1,3'd3,3'd3,3'd2},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1}};

parameter bit [2:0] SpriteTableG_21_35[7:0][7:0] = '{'{3'd3,3'd2,3'd1,3'd3,3'd3,3'd2,3'd0,3'd0},
'{3'd3,3'd1,3'd0,3'd3,3'd3,3'd4,3'd0,3'd0},
'{3'd3,3'd0,3'd0,3'd2,3'd3,3'd0,3'd0,3'd0},
'{3'd3,3'd1,3'd0,3'd4,3'd1,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_22_0[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_22_1[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd3,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_22_2[7:0][7:0] = '{'{3'd0,3'd3,3'd3,3'd2,3'd0,3'd0,3'd4,3'd1},
'{3'd0,3'd3,3'd3,3'd3,3'd2,3'd2,3'd3,3'd3},
'{3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_22_3[7:0][7:0] = '{'{3'd0,3'd2,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2},
'{3'd0,3'd2,3'd3,3'd2,3'd4,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd2,3'd4,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_22_4[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd2,3'd1,3'd0,3'd0,3'd4,3'd1},
'{3'd0,3'd2,3'd2,3'd4,3'd0,3'd0,3'd4,3'd1},
'{3'd2,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd1,3'd4,3'd0,3'd0,3'd0,3'd4},
'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd1,3'd3},
'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd1,3'd3}};

parameter bit [2:0] SpriteTableG_22_5[7:0][7:0] = '{'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd2,3'd4,3'd0,3'd0,3'd0,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd1,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd4,3'd0,3'd3,3'd3},
'{3'd1,3'd2,3'd3,3'd1,3'd0,3'd0,3'd4,3'd1},
'{3'd2,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd0,3'd4,3'd1}};

parameter bit [2:0] SpriteTableG_22_6[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd1,3'd1,3'd3,3'd3},
'{3'd0,3'd2,3'd3,3'd3,3'd4,3'd0,3'd3,3'd1}};

parameter bit [2:0] SpriteTableG_22_7[7:0][7:0] = '{'{3'd1,3'd1,3'd2,3'd4,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd4,3'd1,3'd1,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd3,3'd3},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd1},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd1}};

parameter bit [2:0] SpriteTableG_22_8[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd1},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd0},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd0},
'{3'd2,3'd3,3'd2,3'd2,3'd2,3'd3,3'd3,3'd0},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd1,3'd0},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd1,3'd0},
'{3'd2,3'd3,3'd2,3'd2,3'd3,3'd3,3'd1,3'd0}};

parameter bit [2:0] SpriteTableG_22_9[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd1,3'd2,3'd3,3'd1,3'd0},
'{3'd2,3'd2,3'd2,3'd0,3'd0,3'd3,3'd4,3'd0},
'{3'd2,3'd3,3'd1,3'd0,3'd4,3'd3,3'd4,3'd0},
'{3'd2,3'd3,3'd1,3'd0,3'd1,3'd3,3'd0,3'd0},
'{3'd2,3'd2,3'd1,3'd0,3'd3,3'd3,3'd0,3'd0},
'{3'd2,3'd2,3'd2,3'd2,3'd3,3'd1,3'd0,3'd0},
'{3'd2,3'd3,3'd3,3'd2,3'd3,3'd1,3'd0,3'd0},
'{3'd2,3'd3,3'd2,3'd2,3'd3,3'd1,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_22_10[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd3,3'd1,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd0},
'{3'd3,3'd3,3'd2,3'd3,3'd3,3'd4,3'd0,3'd0},
'{3'd2,3'd3,3'd2,3'd3,3'd3,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_22_11[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd0,3'd0,3'd0,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd0,3'd0,3'd0,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd0,3'd1}};

parameter bit [2:0] SpriteTableG_22_12[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd3},
'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd3},
'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd3},
'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd4,3'd3},
'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd1,3'd3},
'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd1,3'd3},
'{3'd3,3'd3,3'd3,3'd4,3'd0,3'd0,3'd1,3'd3},
'{3'd3,3'd3,3'd3,3'd4,3'd0,3'd0,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_22_13[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd0,3'd0,3'd0,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd0,3'd4,3'd4,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd0,3'd4,3'd1,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd3,3'd3,3'd1,3'd0,3'd1,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd1,3'd0,3'd4,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd1,3'd0,3'd4,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_22_14[7:0][7:0] = '{'{3'd3,3'd3,3'd1,3'd0,3'd1,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd1,3'd0,3'd1,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd4,3'd0,3'd1,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd4,3'd0,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd1,3'd4,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd4,3'd4,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd0,3'd4,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd4,3'd1,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_22_15[7:0][7:0] = '{'{3'd3,3'd3,3'd4,3'd4,3'd2,3'd3,3'd3,3'd3},
'{3'd3,3'd1,3'd0,3'd0,3'd4,3'd3,3'd3,3'd3},
'{3'd3,3'd1,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd1,3'd1,3'd0,3'd2,3'd3,3'd3},
'{3'd3,3'd1,3'd1,3'd1,3'd0,3'd2,3'd3,3'd3},
'{3'd3,3'd1,3'd1,3'd1,3'd0,3'd1,3'd3,3'd3},
'{3'd3,3'd1,3'd3,3'd1,3'd0,3'd4,3'd3,3'd3},
'{3'd3,3'd1,3'd3,3'd3,3'd0,3'd1,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_22_16[7:0][7:0] = '{'{3'd3,3'd4,3'd3,3'd3,3'd0,3'd2,3'd3,3'd3},
'{3'd3,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd1,3'd1,3'd1},
'{3'd0,3'd4,3'd4,3'd0,3'd4,3'd0,3'd0,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_22_17[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3},
'{3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_22_18[7:0][7:0] = '{'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd2,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3},
'{3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_22_19[7:0][7:0] = '{'{3'd1,3'd4,3'd1,3'd1,3'd1,3'd1,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd0,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd4,3'd4,3'd0,3'd1},
'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd3},
'{3'd3,3'd3,3'd1,3'd0,3'd4,3'd0,3'd1,3'd3},
'{3'd3,3'd1,3'd0,3'd0,3'd4,3'd4,3'd3,3'd3},
'{3'd1,3'd0,3'd0,3'd0,3'd4,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_22_20[7:0][7:0] = '{'{3'd0,3'd4,3'd0,3'd4,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd4,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_22_21[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_22_22[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1}};

parameter bit [2:0] SpriteTableG_22_23[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_22_24[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd0,3'd2,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_22_25[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd4,3'd3,3'd3,3'd1,3'd0,3'd4},
'{3'd3,3'd3,3'd4,3'd0,3'd4,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_22_26[7:0][7:0] = '{'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd3},
'{3'd0,3'd0,3'd4,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_22_27[7:0][7:0] = '{'{3'd3,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_22_28[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_22_29[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd1,3'd2,3'd2,3'd2,3'd3,3'd3,3'd1,3'd1},
'{3'd0,3'd2,3'd2,3'd2,3'd3,3'd3,3'd1,3'd1},
'{3'd0,3'd1,3'd2,3'd3,3'd3,3'd2,3'd1,3'd4},
'{3'd0,3'd0,3'd2,3'd3,3'd3,3'd2,3'd1,3'd0}};

parameter bit [2:0] SpriteTableG_22_30[7:0][7:0] = '{'{3'd0,3'd0,3'd1,3'd3,3'd2,3'd2,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd3,3'd2,3'd1,3'd4,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd4,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd3,3'd4,3'd0},
'{3'd1,3'd1,3'd1,3'd4,3'd0,3'd1,3'd4,3'd0},
'{3'd1,3'd1,3'd1,3'd0,3'd0,3'd1,3'd1,3'd0},
'{3'd1,3'd1,3'd1,3'd0,3'd0,3'd4,3'd3,3'd4}};

parameter bit [2:0] SpriteTableG_22_31[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd2,3'd3},
'{3'd0,3'd1,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd3,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_22_32[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd2,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd0,3'd0,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2}};

parameter bit [2:0] SpriteTableG_22_33[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd4,3'd2,3'd3,3'd3,3'd3},
'{3'd0,3'd4,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_22_34[7:0][7:0] = '{'{3'd0,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3},
'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_22_35[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_23_0[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_23_1[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_23_2[7:0][7:0] = '{'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd3},
'{3'd0,3'd0,3'd0,3'd1,3'd2,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd0,3'd1,3'd2,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_23_3[7:0][7:0] = '{'{3'd1,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_23_4[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd4},
'{3'd0,3'd0,3'd0,3'd1,3'd4,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd0,3'd0},
'{3'd0,3'd4,3'd0,3'd4,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd0,3'd4,3'd3,3'd1,3'd0,3'd0,3'd1},
'{3'd4,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd4}};

parameter bit [2:0] SpriteTableG_23_5[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd4,3'd4,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd4,3'd3,3'd3,3'd4,3'd2,3'd3},
'{3'd1,3'd0,3'd4,3'd3,3'd3,3'd4,3'd2,3'd3},
'{3'd0,3'd0,3'd0,3'd1,3'd4,3'd0,3'd0,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2},
'{3'd0,3'd0,3'd0,3'd4,3'd4,3'd0,3'd0,3'd2}};

parameter bit [2:0] SpriteTableG_23_6[7:0][7:0] = '{'{3'd1,3'd0,3'd1,3'd3,3'd3,3'd4,3'd0,3'd3},
'{3'd3,3'd0,3'd1,3'd3,3'd3,3'd1,3'd0,3'd3},
'{3'd2,3'd0,3'd4,3'd3,3'd1,3'd0,3'd0,3'd1},
'{3'd3,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd2,3'd4,3'd1,3'd1,3'd0,3'd0,3'd4},
'{3'd3,3'd0,3'd1,3'd3,3'd3,3'd1,3'd0,3'd3},
'{3'd3,3'd0,3'd1,3'd3,3'd3,3'd1,3'd0,3'd3},
'{3'd1,3'd0,3'd0,3'd1,3'd3,3'd4,3'd0,3'd1}};

parameter bit [2:0] SpriteTableG_23_7[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd4,3'd4,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd4,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd4,3'd1,3'd4,3'd4,3'd4,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd1,3'd1,3'd3}};

parameter bit [2:0] SpriteTableG_23_8[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd2,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd3,3'd3,3'd2,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd3,3'd3,3'd2,3'd2},
'{3'd0,3'd0,3'd0,3'd4,3'd3,3'd3,3'd2,3'd2},
'{3'd0,3'd0,3'd0,3'd1,3'd3,3'd2,3'd2,3'd2},
'{3'd0,3'd0,3'd0,3'd1,3'd3,3'd2,3'd2,3'd2},
'{3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd2,3'd2}};

parameter bit [2:0] SpriteTableG_23_9[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd3,3'd3,3'd2,3'd2,3'd2},
'{3'd0,3'd0,3'd0,3'd3,3'd3,3'd2,3'd2,3'd2},
'{3'd0,3'd0,3'd4,3'd3,3'd3,3'd3,3'd2,3'd2},
'{3'd0,3'd0,3'd1,3'd3,3'd2,3'd3,3'd2,3'd2},
'{3'd0,3'd0,3'd1,3'd3,3'd2,3'd2,3'd2,3'd2},
'{3'd0,3'd0,3'd1,3'd3,3'd2,3'd2,3'd2,3'd2},
'{3'd0,3'd0,3'd3,3'd3,3'd2,3'd3,3'd3,3'd2},
'{3'd0,3'd0,3'd3,3'd3,3'd2,3'd3,3'd2,3'd2}};

parameter bit [2:0] SpriteTableG_23_10[7:0][7:0] = '{'{3'd0,3'd4,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2},
'{3'd0,3'd4,3'd3,3'd3,3'd2,3'd3,3'd3,3'd2},
'{3'd0,3'd1,3'd3,3'd3,3'd2,3'd3,3'd3,3'd2},
'{3'd0,3'd1,3'd3,3'd2,3'd2,3'd3,3'd2,3'd3},
'{3'd0,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd2},
'{3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_23_11[7:0][7:0] = '{'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_23_12[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_23_13[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_23_14[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_23_15[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_23_16[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd1,3'd1,3'd1,3'd4,3'd0,3'd0},
'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd3}};

parameter bit [2:0] SpriteTableG_23_17[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd1,3'd1,3'd1,3'd4,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd0,3'd0},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd3,3'd3,3'd2,3'd2,3'd3,3'd3,3'd3},
'{3'd2,3'd3,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_23_18[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd3,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd3,3'd3,3'd2,3'd1,3'd3,3'd3,3'd3},
'{3'd2,3'd3,3'd3,3'd1,3'd0,3'd1,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd2,3'd0,3'd0,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_23_19[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_23_20[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd0},
'{3'd3,3'd3,3'd3,3'd1,3'd3,3'd1,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_23_21[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd0,3'd1},
'{3'd3,3'd0,3'd4,3'd4,3'd0,3'd0,3'd4,3'd3},
'{3'd3,3'd4,3'd0,3'd0,3'd0,3'd0,3'd3,3'd3},
'{3'd3,3'd1,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd1,3'd0,3'd4,3'd0,3'd1,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_23_22[7:0][7:0] = '{'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_23_23[7:0][7:0] = '{'{3'd0,3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd0,3'd0,3'd0,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd1,3'd4,3'd0,3'd1,3'd3,3'd3,3'd3},
'{3'd3,3'd1,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd0,3'd0,3'd0,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd1,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_23_24[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd4,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd1,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd0,3'd4,3'd4,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd0,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd1,3'd0}};

parameter bit [2:0] SpriteTableG_23_25[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd1,3'd4,3'd0},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd1,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd1,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_23_26[7:0][7:0] = '{'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd1,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd4,3'd0,3'd0},
'{3'd3,3'd3,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0},
'{3'd3,3'd1,3'd2,3'd3,3'd3,3'd4,3'd0,3'd1},
'{3'd3,3'd2,3'd3,3'd3,3'd3,3'd1,3'd0,3'd3},
'{3'd3,3'd3,3'd2,3'd3,3'd3,3'd4,3'd0,3'd1}};

parameter bit [2:0] SpriteTableG_23_27[7:0][7:0] = '{'{3'd3,3'd3,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd1,3'd1,3'd1,3'd0,3'd0,3'd4},
'{3'd3,3'd3,3'd2,3'd3,3'd3,3'd4,3'd0,3'd1},
'{3'd3,3'd3,3'd1,3'd0,3'd4,3'd0,3'd0,3'd1},
'{3'd3,3'd3,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd2,3'd4,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_23_28[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd0,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd0,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd0,3'd0},
'{3'd3,3'd3,3'd2,3'd2,3'd1,3'd4,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_23_29[7:0][7:0] = '{'{3'd1,3'd0,3'd1,3'd4,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_23_30[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_23_31[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd1,3'd4,3'd0,3'd0,3'd4,3'd4,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd4,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd3,3'd3,3'd2,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd3,3'd3,3'd2,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_23_32[7:0][7:0] = '{'{3'd2,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd3,3'd3,3'd4,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd3,3'd4,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd2,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd2,3'd3,3'd4,3'd0,3'd0,3'd0},
'{3'd2,3'd3,3'd2,3'd2,3'd3,3'd4,3'd0,3'd0},
'{3'd2,3'd3,3'd3,3'd2,3'd2,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_23_33[7:0][7:0] = '{'{3'd2,3'd3,3'd3,3'd3,3'd2,3'd2,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_23_34[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_23_35[7:0][7:0] = '{'{3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd0,3'd2,3'd3,3'd3,3'd3,3'd3,3'd2,3'd0},
'{3'd0,3'd2,3'd3,3'd3,3'd3,3'd3,3'd0,3'd0},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0},
'{3'd0,3'd1,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd4,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd4,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_24_0[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd2,3'd3,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd2,3'd3,3'd2,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_24_1[7:0][7:0] = '{'{3'd0,3'd0,3'd2,3'd3,3'd3,3'd2,3'd0,3'd0},
'{3'd0,3'd0,3'd3,3'd3,3'd3,3'd3,3'd2,3'd0},
'{3'd0,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_24_2[7:0][7:0] = '{'{3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd0,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_24_3[7:0][7:0] = '{'{3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_24_4[7:0][7:0] = '{'{3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4},
'{3'd4,3'd0,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd0,3'd0,3'd2,3'd3,3'd3,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd2,3'd3,3'd2,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd4,3'd4,3'd0,3'd1,3'd1,3'd0,3'd0},
'{3'd3,3'd4,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_24_5[7:0][7:0] = '{'{3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd3,3'd2,3'd4,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd2,3'd4,3'd4,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd1,3'd2,3'd3,3'd4,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_24_6[7:0][7:0] = '{'{3'd3,3'd1,3'd0,3'd1,3'd3,3'd3,3'd0,3'd0},
'{3'd3,3'd1,3'd0,3'd4,3'd3,3'd3,3'd4,3'd0},
'{3'd3,3'd4,3'd0,3'd0,3'd1,3'd2,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd4,3'd4,3'd0,3'd1},
'{3'd3,3'd1,3'd0,3'd4,3'd3,3'd3,3'd1,3'd1},
'{3'd3,3'd3,3'd0,3'd1,3'd3,3'd3,3'd1,3'd0},
'{3'd3,3'd1,3'd0,3'd0,3'd1,3'd3,3'd4,3'd0}};

parameter bit [2:0] SpriteTableG_24_7[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd1,3'd4,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0},
'{3'd3,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd4,3'd4,3'd4,3'd1,3'd1,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_24_8[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd3,3'd2,3'd2,3'd3,3'd2,3'd2,3'd3,3'd2}};

parameter bit [2:0] SpriteTableG_24_9[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd3,3'd2,3'd2,3'd3,3'd2,3'd2,3'd3,3'd2},
'{3'd3,3'd2,3'd2,3'd3,3'd2,3'd2,3'd3,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3},
'{3'd3,3'd3,3'd2,3'd3,3'd3,3'd2,3'd3,3'd3},
'{3'd2,3'd2,3'd2,3'd2,3'd3,3'd2,3'd2,3'd3}};

parameter bit [2:0] SpriteTableG_24_10[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd3,3'd2,3'd2,3'd2,3'd3,3'd2,3'd2,3'd3},
'{3'd3,3'd3,3'd2,3'd3,3'd2,3'd2,3'd2,3'd3},
'{3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3},
'{3'd3,3'd2,3'd2,3'd2,3'd3,3'd2,3'd2,3'd1},
'{3'd3,3'd3,3'd2,3'd2,3'd3,3'd2,3'd3,3'd1},
'{3'd3,3'd2,3'd2,3'd2,3'd3,3'd2,3'd3,3'd1},
'{3'd3,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd1}};

parameter bit [2:0] SpriteTableG_24_11[7:0][7:0] = '{'{3'd3,3'd3,3'd2,3'd2,3'd3,3'd2,3'd3,3'd1},
'{3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd3,3'd4},
'{3'd3,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3},
'{3'd3,3'd3,3'd2,3'd3,3'd3,3'd2,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_24_12[7:0][7:0] = '{'{3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd2,3'd2,3'd3,3'd2,3'd2,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_24_13[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd0,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd0,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd0,3'd3}};

parameter bit [2:0] SpriteTableG_24_14[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd4,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd1,3'd3},
'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd1,3'd1},
'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd1,3'd4,3'd0,3'd1,3'd4},
'{3'd3,3'd3,3'd3,3'd4,3'd0,3'd0,3'd0,3'd4},
'{3'd3,3'd3,3'd3,3'd1,3'd1,3'd1,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_24_15[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_24_16[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd4,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd1},
'{3'd4,3'd1,3'd1,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_24_17[7:0][7:0] = '{'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd1,3'd1,3'd1,3'd4},
'{3'd0,3'd0,3'd1,3'd3,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd3,3'd3,3'd3,3'd0,3'd0},
'{3'd4,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd0},
'{3'd3,3'd0,3'd0,3'd0,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd1,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd0,3'd0,3'd4,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_24_18[7:0][7:0] = '{'{3'd3,3'd3,3'd4,3'd0,3'd0,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd1,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_24_19[7:0][7:0] = '{'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd4,3'd0,3'd0,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd0,3'd0,3'd4,3'd3,3'd3,3'd3},
'{3'd3,3'd1,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3},
'{3'd3,3'd1,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3},
'{3'd3,3'd0,3'd0,3'd0,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_24_20[7:0][7:0] = '{'{3'd1,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd0,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_24_21[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd1,3'd1,3'd3},
'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd1,3'd1,3'd4},
'{3'd3,3'd3,3'd3,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd3,3'd3,3'd1,3'd4,3'd4,3'd0,3'd0,3'd4},
'{3'd3,3'd3,3'd3,3'd1,3'd1,3'd4,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_24_22[7:0][7:0] = '{'{3'd3,3'd2,3'd0,3'd1,3'd1,3'd1,3'd4,3'd0},
'{3'd1,3'd0,3'd1,3'd0,3'd2,3'd4,3'd1,3'd4},
'{3'd0,3'd0,3'd1,3'd0,3'd0,3'd2,3'd4,3'd1},
'{3'd0,3'd1,3'd0,3'd0,3'd1,3'd0,3'd2,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd0,3'd1,3'd0,3'd2},
'{3'd2,3'd0,3'd1,3'd0,3'd1,3'd0,3'd1,3'd1},
'{3'd3,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_24_23[7:0][7:0] = '{'{3'd3,3'd3,3'd0,3'd1,3'd0,3'd0,3'd0,3'd1},
'{3'd3,3'd3,3'd2,3'd0,3'd0,3'd1,3'd0,3'd1},
'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd0,3'd0,3'd0,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd0,3'd0,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0},
'{3'd3,3'd2,3'd3,3'd3,3'd3,3'd2,3'd0,3'd0},
'{3'd3,3'd2,3'd0,3'd1,3'd2,3'd3,3'd1,3'd0}};

parameter bit [2:0] SpriteTableG_24_24[7:0][7:0] = '{'{3'd3,3'd3,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0},
'{3'd3,3'd3,3'd2,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd3,3'd3,3'd3,3'd0,3'd1,3'd0,3'd0,3'd1},
'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd1,3'd1,3'd1},
'{3'd3,3'd3,3'd1,3'd1,3'd0,3'd1,3'd1,3'd1},
'{3'd3,3'd3,3'd3,3'd2,3'd1,3'd1,3'd1,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd1,3'd1,3'd0},
'{3'd1,3'd3,3'd1,3'd3,3'd2,3'd1,3'd1,3'd1}};

parameter bit [2:0] SpriteTableG_24_25[7:0][7:0] = '{'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd1,3'd1,3'd1},
'{3'd0,3'd3,3'd3,3'd3,3'd3,3'd1,3'd1,3'd1},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd2,3'd0,3'd0},
'{3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd1,3'd2,3'd2},
'{3'd1,3'd4,3'd1,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_24_26[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd0,3'd1,3'd3,3'd3,3'd2,3'd0},
'{3'd3,3'd1,3'd0,3'd4,3'd1,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd1,3'd0,3'd4,3'd3,3'd1,3'd0,3'd0},
'{3'd3,3'd1,3'd0,3'd4,3'd3,3'd3,3'd4,3'd0},
'{3'd3,3'd4,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_24_27[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd4,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0},
'{3'd3,3'd1,3'd0,3'd0,3'd3,3'd3,3'd0,3'd0},
'{3'd3,3'd4,3'd0,3'd0,3'd2,3'd2,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd2},
'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2},
'{3'd4,3'd0,3'd0,3'd1,3'd1,3'd1,3'd2,3'd1}};

parameter bit [2:0] SpriteTableG_24_28[7:0][7:0] = '{'{3'd3,3'd4,3'd0,3'd1,3'd3,3'd3,3'd1,3'd1},
'{3'd1,3'd0,3'd0,3'd2,3'd3,3'd3,3'd2,3'd2},
'{3'd4,3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_24_29[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_24_30[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_24_31[7:0][7:0] = '{'{3'd0,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_24_32[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd4,3'd0,3'd0},
'{3'd4,3'd0,3'd0,3'd0,3'd4,3'd4,3'd0,3'd0},
'{3'd1,3'd4,3'd0,3'd4,3'd4,3'd0,3'd0,3'd0},
'{3'd4,3'd1,3'd1,3'd4,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_24_33[7:0][7:0] = '{'{3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd4,3'd2},
'{3'd3,3'd3,3'd1,3'd4,3'd1,3'd2,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_24_34[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_24_35[7:0][7:0] = '{'{3'd2,3'd0,3'd0,3'd4,3'd1,3'd1,3'd2,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_25_0[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_25_1[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd1,3'd0,3'd0,3'd4,3'd1,3'd2,3'd2},
'{3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_25_2[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_25_3[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd2,3'd1,3'd2,3'd2,3'd3,3'd3,3'd3},
'{3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd1}};

parameter bit [2:0] SpriteTableG_25_4[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd1,3'd0,3'd0,3'd0,3'd4,3'd4,3'd0},
'{3'd0,3'd1,3'd0,3'd0,3'd0,3'd4,3'd4,3'd0}};

parameter bit [2:0] SpriteTableG_25_5[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd1},
'{3'd4,3'd3,3'd4,3'd0,3'd0,3'd2,3'd3,3'd2},
'{3'd1,3'd3,3'd4,3'd0,3'd0,3'd3,3'd3,3'd2},
'{3'd0,3'd4,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1}};

parameter bit [2:0] SpriteTableG_25_6[7:0][7:0] = '{'{3'd1,3'd3,3'd1,3'd0,3'd1,3'd3,3'd3,3'd1},
'{3'd1,3'd3,3'd1,3'd0,3'd1,3'd3,3'd3,3'd1},
'{3'd4,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd1},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd2,3'd3,3'd2,3'd1,3'd1,3'd3,3'd2,3'd1},
'{3'd3,3'd3,3'd3,3'd1,3'd1,3'd2,3'd1,3'd0},
'{3'd1,3'd3,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_25_7[7:0][7:0] = '{'{3'd1,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd1,3'd1},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2}};

parameter bit [2:0] SpriteTableG_25_8[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableG_25_9[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd4,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1},
'{3'd3,3'd4,3'd0,3'd4,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd0,3'd0,3'd4,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_25_10[7:0][7:0] = '{'{3'd1,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd0,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd4,3'd3,3'd3,3'd1,3'd1,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_25_11[7:0][7:0] = '{'{3'd0,3'd4,3'd4,3'd0,3'd4,3'd4,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd0,3'd4},
'{3'd1,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd2,3'd3,3'd2,3'd3,3'd2,3'd2,3'd2},
'{3'd3,3'd3,3'd3,3'd2,3'd3,3'd3,3'd2,3'd3}};

parameter bit [2:0] SpriteTableG_25_12[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd2,3'd3,3'd3,3'd2,3'd2},
'{3'd3,3'd3,3'd2,3'd3,3'd3,3'd2,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd4,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_25_13[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd4,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_25_14[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd4,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd4,3'd4,3'd0,3'd4,3'd4,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd3,3'd3,3'd3,3'd3,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4}};

parameter bit [2:0] SpriteTableG_25_15[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0}};

parameter bit [2:0] SpriteTableG_25_16[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd1,3'd1,3'd1,3'd4,3'd0},
'{3'd4,3'd1,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd4,3'd4,3'd1,3'd1,3'd3},
'{3'd1,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1}};

parameter bit [2:0] SpriteTableG_25_17[7:0][7:0] = '{'{3'd0,3'd4,3'd1,3'd1,3'd4,3'd4,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3},
'{3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3}};

parameter bit [2:0] SpriteTableG_25_18[7:0][7:0] = '{'{3'd3,3'd4,3'd0,3'd0,3'd0,3'd4,3'd3,3'd3},
'{3'd3,3'd1,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd3,3'd3,3'd0,3'd0,3'd0,3'd3,3'd3,3'd1},
'{3'd3,3'd3,3'd4,3'd0,3'd4,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd4,3'd0,3'd1,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd1,3'd0,3'd4,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_25_19[7:0][7:0] = '{'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd3,3'd3},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd1,3'd3},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd3,3'd3,3'd4,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd3,3'd3,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_25_20[7:0][7:0] = '{'{3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd4,3'd1,3'd4,3'd4,3'd4,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_25_21[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd1,3'd4,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd1,3'd1,3'd4,3'd1,3'd2,3'd1,3'd0}};

parameter bit [2:0] SpriteTableG_25_22[7:0][7:0] = '{'{3'd0,3'd4,3'd1,3'd1,3'd4,3'd4,3'd2,3'd2},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd4,3'd1},
'{3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd4},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd2,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd4},
'{3'd3,3'd1,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd1,3'd0,3'd1,3'd1,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_25_23[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd4,3'd0,3'd1,3'd1,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd4,3'd0,3'd1,3'd1},
'{3'd4,3'd1,3'd0,3'd4,3'd1,3'd0,3'd0,3'd1},
'{3'd3,3'd3,3'd3,3'd0,3'd1,3'd3,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd4,3'd1,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd1},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_25_24[7:0][7:0] = '{'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd1,3'd1,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd1,3'd1,3'd1,3'd0,3'd1,3'd3,3'd1,3'd0},
'{3'd1,3'd0,3'd0,3'd1,3'd1,3'd3,3'd4,3'd0},
'{3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_25_25[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd3,3'd2,3'd2,3'd1,3'd0,3'd1,3'd0,3'd0},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd2,3'd0,3'd0},
'{3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd1,3'd1}};

parameter bit [2:0] SpriteTableG_25_26[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd2,3'd0,3'd1,3'd1,3'd1},
'{3'd1,3'd3,3'd3,3'd2,3'd0,3'd3,3'd3,3'd0},
'{3'd4,3'd2,3'd3,3'd1,3'd0,3'd4,3'd4,3'd0},
'{3'd0,3'd0,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd4,3'd4,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd1,3'd4,3'd0,3'd0,3'd1,3'd4,3'd0},
'{3'd1,3'd3,3'd1,3'd0,3'd0,3'd3,3'd3,3'd1},
'{3'd4,3'd1,3'd0,3'd0,3'd1,3'd3,3'd1,3'd1}};

parameter bit [2:0] SpriteTableG_25_27[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd4,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd3,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd2,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_25_28[7:0][7:0] = '{'{3'd1,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd1,3'd4,3'd1,3'd4,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1}};

parameter bit [2:0] SpriteTableG_25_29[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_25_30[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_25_31[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_25_32[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_25_33[7:0][7:0] = '{'{3'd2,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd2,3'd4,3'd0,3'd0,3'd4,3'd1},
'{3'd1,3'd1,3'd2,3'd2,3'd2,3'd3,3'd3,3'd2},
'{3'd1,3'd1,3'd1,3'd1,3'd2,3'd2,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1,3'd1},
'{3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1}};

parameter bit [2:0] SpriteTableG_25_34[7:0][7:0] = '{'{3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd3,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd3,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd3,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0},
'{3'd3,3'd3,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd3,3'd3,3'd2,3'd1,3'd1,3'd1,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_25_35[7:0][7:0] = '{'{3'd3,3'd3,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd4,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_26_0[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_26_1[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd4,3'd1,3'd1,3'd0,3'd0,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd2,3'd0,3'd1,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd2,3'd1,3'd1,3'd1,3'd0},
'{3'd3,3'd3,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd3,3'd3,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1}};

parameter bit [2:0] SpriteTableG_26_2[7:0][7:0] = '{'{3'd3,3'd2,3'd4,3'd2,3'd1,3'd1,3'd1,3'd1},
'{3'd3,3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd0},
'{3'd2,3'd0,3'd4,3'd0,3'd0,3'd1,3'd1,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_26_3[7:0][7:0] = '{'{3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd2,3'd3,3'd2,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_26_4[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd4,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_26_5[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd1,3'd1,3'd4,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd2,3'd2},
'{3'd2,3'd1,3'd1,3'd1,3'd2,3'd2,3'd1,3'd2}};

parameter bit [2:0] SpriteTableG_26_6[7:0][7:0] = '{'{3'd1,3'd2,3'd3,3'd1,3'd1,3'd1,3'd2,3'd2},
'{3'd1,3'd2,3'd3,3'd2,3'd1,3'd1,3'd2,3'd2},
'{3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1},
'{3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd2},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd3},
'{3'd0,3'd0,3'd0,3'd1,3'd0,3'd1,3'd3,3'd3},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2}};

parameter bit [2:0] SpriteTableG_26_7[7:0][7:0] = '{'{3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4},
'{3'd1,3'd1,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3}};

parameter bit [2:0] SpriteTableG_26_8[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd1},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd1},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd4},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd0},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd0}};

parameter bit [2:0] SpriteTableG_26_9[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd3,3'd2,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd4,3'd4,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_26_10[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd4,3'd1,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1},
'{3'd2,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd0,3'd1,3'd1,3'd1,3'd0,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2}};

parameter bit [2:0] SpriteTableG_26_11[7:0][7:0] = '{'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd4,3'd4,3'd4,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd1,3'd3,3'd1,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd3,3'd3,3'd1,3'd4,3'd0,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd4,3'd0,3'd0,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd4,3'd0,3'd4,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd4,3'd4,3'd4,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_26_12[7:0][7:0] = '{'{3'd3,3'd1,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3},
'{3'd3,3'd1,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3},
'{3'd3,3'd1,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3},
'{3'd3,3'd1,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3},
'{3'd3,3'd1,3'd0,3'd0,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd4,3'd0,3'd0,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd0,3'd0,3'd4,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd4,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_26_13[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd4,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd1,3'd4},
'{3'd0,3'd0,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0}};

parameter bit [2:0] SpriteTableG_26_14[7:0][7:0] = '{'{3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd0},
'{3'd0,3'd0,3'd3,3'd3,3'd3,3'd3,3'd2,3'd0},
'{3'd0,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd4,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd0,3'd0,3'd0,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1}};

parameter bit [2:0] SpriteTableG_26_15[7:0][7:0] = '{'{3'd4,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd1,3'd1},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0}};

parameter bit [2:0] SpriteTableG_26_16[7:0][7:0] = '{'{3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd0},
'{3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd0},
'{3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0},
'{3'd1,3'd1,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_26_17[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd1,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_26_18[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd0,3'd1},
'{3'd3,3'd3,3'd3,3'd2,3'd1,3'd1,3'd0,3'd1},
'{3'd3,3'd3,3'd2,3'd0,3'd1,3'd1,3'd1,3'd0},
'{3'd3,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_26_19[7:0][7:0] = '{'{3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd1,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd1},
'{3'd0,3'd4,3'd3,3'd3,3'd3,3'd1,3'd1,3'd0},
'{3'd0,3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd1}};

parameter bit [2:0] SpriteTableG_26_20[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd4,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd3,3'd1,3'd1,3'd1,3'd1,3'd4,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_26_21[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd1,3'd2,3'd2,3'd2,3'd3}};

parameter bit [2:0] SpriteTableG_26_22[7:0][7:0] = '{'{3'd1,3'd1,3'd2,3'd1,3'd0,3'd0,3'd1,3'd2},
'{3'd1,3'd3,3'd3,3'd3,3'd0,3'd4,3'd3,3'd3},
'{3'd4,3'd3,3'd3,3'd3,3'd0,3'd1,3'd3,3'd3},
'{3'd1,3'd0,3'd1,3'd3,3'd1,3'd1,3'd3,3'd3},
'{3'd1,3'd1,3'd0,3'd4,3'd3,3'd2,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd4,3'd0,3'd1,3'd3,3'd2},
'{3'd4,3'd1,3'd1,3'd1,3'd1,3'd0,3'd1,3'd3},
'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd4}};

parameter bit [2:0] SpriteTableG_26_23[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd1,3'd3},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd3,3'd3,3'd0},
'{3'd0,3'd1,3'd1,3'd0,3'd1,3'd3,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd1,3'd3,3'd4,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd1,3'd3,3'd0,3'd0,3'd0},
'{3'd3,3'd4,3'd0,3'd3,3'd1,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_26_24[7:0][7:0] = '{'{3'd3,3'd3,3'd4,3'd3,3'd4,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd4,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd1,3'd1,3'd1,3'd1,3'd0},
'{3'd1,3'd4,3'd0,3'd0,3'd0,3'd0,3'd4,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_26_25[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_26_26[7:0][7:0] = '{'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd1,3'd1,3'd1,3'd4,3'd4,3'd1,3'd1,3'd1},
'{3'd0,3'd4,3'd1,3'd1,3'd1,3'd3,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd2,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd3,3'd3,3'd2},
'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd3,3'd3,3'd3},
'{3'd1,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd4,3'd0,3'd0,3'd4,3'd1,3'd2,3'd3}};

parameter bit [2:0] SpriteTableG_26_27[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd4,3'd4},
'{3'd0,3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_26_28[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd4,3'd4,3'd1,3'd1,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_26_29[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_26_30[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_26_31[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_26_32[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd0,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd4,3'd0,3'd4,3'd2,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd2,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd4,3'd2,3'd1,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_26_33[7:0][7:0] = '{'{3'd0,3'd0,3'd1,3'd2,3'd1,3'd1,3'd0,3'd0},
'{3'd4,3'd1,3'd2,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd3,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0},
'{3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1,3'd0},
'{3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1}};

parameter bit [2:0] SpriteTableG_26_34[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_26_35[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_27_0[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_27_1[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_27_2[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd0,3'd0,3'd4}};

parameter bit [2:0] SpriteTableG_27_3[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd2,3'd2,3'd1,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd2,3'd3,3'd3,3'd3},
'{3'd0,3'd4,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3},
'{3'd0,3'd2,3'd1,3'd0,3'd1,3'd3,3'd3,3'd3},
'{3'd0,3'd2,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd2,3'd3,3'd3,3'd3,3'd1,3'd2,3'd3},
'{3'd0,3'd2,3'd3,3'd3,3'd3,3'd2,3'd2,3'd3},
'{3'd0,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_27_4[7:0][7:0] = '{'{3'd0,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_27_5[7:0][7:0] = '{'{3'd0,3'd0,3'd2,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd0,3'd0,3'd2,3'd3,3'd3,3'd3,3'd2,3'd0},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd3,3'd3,3'd1,3'd1,3'd2},
'{3'd0,3'd0,3'd0,3'd3,3'd2,3'd0,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd4,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd1,3'd0,3'd0,3'd0,3'd1,3'd2,3'd0}};

parameter bit [2:0] SpriteTableG_27_6[7:0][7:0] = '{'{3'd2,3'd2,3'd1,3'd4,3'd2,3'd3,3'd3,3'd0},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd1}};

parameter bit [2:0] SpriteTableG_27_7[7:0][7:0] = '{'{3'd1,3'd1,3'd3,3'd3,3'd2,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd1,3'd1,3'd0,3'd0,3'd4,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd1,3'd3},
'{3'd4,3'd0,3'd0,3'd0,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd0,3'd0,3'd4,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_27_8[7:0][7:0] = '{'{3'd4,3'd0,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd4,3'd3,3'd3,3'd1,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd1,3'd3,3'd3,3'd2}};

parameter bit [2:0] SpriteTableG_27_9[7:0][7:0] = '{'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_27_10[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd2,3'd3,3'd3,3'd1,3'd3},
'{3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2,3'd2},
'{3'd0,3'd0,3'd1,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_27_11[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd1},
'{3'd3,3'd3,3'd3,3'd1,3'd4,3'd4,3'd0,3'd0},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd3},
'{3'd3,3'd3,3'd4,3'd0,3'd0,3'd0,3'd1,3'd3},
'{3'd3,3'd3,3'd4,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd3,3'd3,3'd4,3'd0,3'd1,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_27_12[7:0][7:0] = '{'{3'd3,3'd3,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd1,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd1,3'd1,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0}};

parameter bit [2:0] SpriteTableG_27_13[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd2,3'd0,3'd0,3'd1,3'd1},
'{3'd3,3'd3,3'd3,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd3,3'd3,3'd1,3'd1,3'd0,3'd1,3'd0,3'd0},
'{3'd3,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1},
'{3'd2,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd1,3'd0,3'd1,3'd1,3'd1,3'd0,3'd1,3'd0}};

parameter bit [2:0] SpriteTableG_27_14[7:0][7:0] = '{'{3'd0,3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd1,3'd1},
'{3'd1,3'd0,3'd1,3'd0,3'd0,3'd1,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd0,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_27_15[7:0][7:0] = '{'{3'd1,3'd1,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0},
'{3'd3,3'd2,3'd1,3'd0,3'd0,3'd1,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd2,3'd1,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd0},
'{3'd4,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_27_16[7:0][7:0] = '{'{3'd0,3'd0,3'd4,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd1,3'd3,3'd3},
'{3'd0,3'd0,3'd4,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_27_17[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd0}};

parameter bit [2:0] SpriteTableG_27_18[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd2,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd2,3'd0,3'd0,3'd1,3'd0,3'd0,3'd1},
'{3'd1,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0},
'{3'd1,3'd0,3'd1,3'd1,3'd0,3'd1,3'd0,3'd2},
'{3'd1,3'd0,3'd1,3'd1,3'd0,3'd0,3'd1,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd1,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd3}};

parameter bit [2:0] SpriteTableG_27_19[7:0][7:0] = '{'{3'd0,3'd1,3'd1,3'd0,3'd1,3'd0,3'd4,3'd3},
'{3'd0,3'd1,3'd1,3'd0,3'd1,3'd0,3'd1,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd3,3'd3},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd4,3'd4,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd1,3'd0,3'd3},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd1,3'd0,3'd1},
'{3'd0,3'd1,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_27_20[7:0][7:0] = '{'{3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0},
'{3'd3,3'd3,3'd1,3'd0,3'd1,3'd1,3'd1,3'd1},
'{3'd3,3'd3,3'd3,3'd2,3'd0,3'd0,3'd0,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd2,3'd0},
'{3'd1,3'd1,3'd1,3'd3,3'd1,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0}};

parameter bit [2:0] SpriteTableG_27_21[7:0][7:0] = '{'{3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd0,3'd0,3'd1,3'd1,3'd2,3'd3,3'd3},
'{3'd3,3'd3,3'd1,3'd0,3'd1,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd2,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_27_22[7:0][7:0] = '{'{3'd1,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd1,3'd2,3'd3,3'd3,3'd3,3'd1,3'd4},
'{3'd2,3'd1,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd3,3'd1,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd2,3'd3,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd2,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd3,3'd3,3'd4,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_27_23[7:0][7:0] = '{'{3'd1,3'd3,3'd3,3'd4,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd1,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd4,3'd4,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_27_24[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_27_25[7:0][7:0] = '{'{3'd0,3'd0,3'd4,3'd4,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd4,3'd4,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd4,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd4,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd3,3'd1,3'd3,3'd1,3'd1,3'd1},
'{3'd4,3'd3,3'd4,3'd0,3'd1,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_27_26[7:0][7:0] = '{'{3'd3,3'd1,3'd0,3'd1,3'd2,3'd1,3'd1,3'd1},
'{3'd4,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd1,3'd1,3'd1},
'{3'd0,3'd4,3'd1,3'd2,3'd1,3'd1,3'd0,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd2,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd2,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_27_27[7:0][7:0] = '{'{3'd1,3'd2,3'd2,3'd0,3'd0,3'd0,3'd4,3'd1},
'{3'd1,3'd1,3'd3,3'd2,3'd2,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd4,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_27_28[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_27_29[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd4,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_27_30[7:0][7:0] = '{'{3'd0,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd4,3'd1,3'd4,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_27_31[7:0][7:0] = '{'{3'd0,3'd4,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd4,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd1,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd1,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_27_32[7:0][7:0] = '{'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd1,3'd1,3'd1,3'd4,3'd4,3'd1,3'd1},
'{3'd0,3'd0,3'd4,3'd4,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_27_33[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3}};

parameter bit [2:0] SpriteTableG_27_34[7:0][7:0] = '{'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_27_35[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_28_0[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_28_1[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1}};

parameter bit [2:0] SpriteTableG_28_2[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd4,3'd3,3'd3,3'd1,3'd1},
'{3'd0,3'd0,3'd4,3'd3,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd3,3'd4,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd4,3'd3,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd2,3'd3,3'd0,3'd0,3'd0,3'd0,3'd1,3'd4}};

parameter bit [2:0] SpriteTableG_28_3[7:0][7:0] = '{'{3'd3,3'd3,3'd4,3'd0,3'd0,3'd0,3'd1,3'd4},
'{3'd3,3'd1,3'd1,3'd0,3'd0,3'd0,3'd4,3'd1},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd3,3'd3,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd1,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_28_4[7:0][7:0] = '{'{3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd4,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3},
'{3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd4,3'd1},
'{3'd3,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd2,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd2,3'd2,3'd2,3'd0,3'd0,3'd1,3'd1},
'{3'd3,3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1}};

parameter bit [2:0] SpriteTableG_28_5[7:0][7:0] = '{'{3'd1,3'd2,3'd2,3'd2,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0},
'{3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_28_6[7:0][7:0] = '{'{3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3},
'{3'd1,3'd0,3'd0,3'd0,3'd4,3'd2,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_28_7[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2},
'{3'd2,3'd1,3'd0,3'd0,3'd1,3'd2,3'd1,3'd1},
'{3'd3,3'd3,3'd1,3'd1,3'd3,3'd2,3'd1,3'd1},
'{3'd3,3'd3,3'd1,3'd2,3'd2,3'd1,3'd1,3'd1},
'{3'd3,3'd2,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd3,3'd2,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd3,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_28_8[7:0][7:0] = '{'{3'd3,3'd1,3'd1,3'd1,3'd3,3'd2,3'd0,3'd0},
'{3'd3,3'd1,3'd1,3'd1,3'd2,3'd1,3'd1,3'd0},
'{3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd0,3'd0,3'd4,3'd3,3'd1,3'd0,3'd0},
'{3'd2,3'd1,3'd0,3'd4,3'd3,3'd4,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_28_9[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd0,3'd4,3'd2,3'd1},
'{3'd2,3'd2,3'd2,3'd0,3'd0,3'd0,3'd2,3'd3},
'{3'd3,3'd2,3'd1,3'd4,3'd3,3'd2,3'd2,3'd3},
'{3'd3,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd3,3'd3,3'd2,3'd0},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd1,3'd1},
'{3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd0,3'd2},
'{3'd3,3'd2,3'd2,3'd3,3'd3,3'd2,3'd0,3'd3}};

parameter bit [2:0] SpriteTableG_28_10[7:0][7:0] = '{'{3'd3,3'd3,3'd2,3'd3,3'd3,3'd1,3'd4,3'd2},
'{3'd3,3'd3,3'd2,3'd2,3'd3,3'd2,3'd1,3'd0},
'{3'd2,3'd2,3'd1,3'd1,3'd1,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd1,3'd1,3'd2,3'd2,3'd2,3'd3},
'{3'd1,3'd2,3'd2,3'd2,3'd3,3'd3,3'd1,3'd1},
'{3'd3,3'd3,3'd0,3'd0,3'd4,3'd1,3'd3,3'd3},
'{3'd3,3'd3,3'd1,3'd1,3'd1,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd1,3'd4,3'd1,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_28_11[7:0][7:0] = '{'{3'd4,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd4,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd4,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd1,3'd4,3'd1,3'd3,3'd3,3'd3,3'd1,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd1,3'd1}};

parameter bit [2:0] SpriteTableG_28_12[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd1,3'd1,3'd1},
'{3'd3,3'd3,3'd3,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd2,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_28_13[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0},
'{3'd0,3'd1,3'd0,3'd1,3'd2,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd1,3'd1,3'd4,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd0,3'd4,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd1,3'd3,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd4,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_28_14[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd4,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd4,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0},
'{3'd0,3'd1,3'd1,3'd2,3'd3,3'd2,3'd1,3'd0},
'{3'd1,3'd1,3'd1,3'd3,3'd3,3'd2,3'd0,3'd0},
'{3'd1,3'd0,3'd1,3'd2,3'd3,3'd4,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_28_15[7:0][7:0] = '{'{3'd0,3'd1,3'd0,3'd0,3'd3,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd2,3'd3,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0},
'{3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd1},
'{3'd3,3'd2,3'd1,3'd0,3'd0,3'd1,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_28_16[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd0}};

parameter bit [2:0] SpriteTableG_28_17[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd0,3'd0},
'{3'd3,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_28_18[7:0][7:0] = '{'{3'd0,3'd1,3'd1,3'd1,3'd2,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd1,3'd2,3'd0,3'd0,3'd1},
'{3'd0,3'd1,3'd0,3'd0,3'd0,3'd4,3'd1,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd3,3'd2,3'd1,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd1,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2}};

parameter bit [2:0] SpriteTableG_28_19[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd2,3'd3,3'd3,3'd1,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd1},
'{3'd2,3'd2,3'd3,3'd3,3'd3,3'd4,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd4,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd2,3'd3,3'd0,3'd0,3'd0},
'{3'd3,3'd4,3'd0,3'd4,3'd3,3'd1,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd1,3'd4,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_28_20[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0},
'{3'd3,3'd4,3'd0,3'd4,3'd3,3'd3,3'd1,3'd0},
'{3'd2,3'd0,3'd0,3'd0,3'd3,3'd3,3'd3,3'd1},
'{3'd0,3'd1,3'd0,3'd0,3'd2,3'd2,3'd2,3'd2},
'{3'd1,3'd0,3'd1,3'd0,3'd2,3'd2,3'd2,3'd2},
'{3'd3,3'd2,3'd1,3'd0,3'd2,3'd3,3'd3,3'd2},
'{3'd3,3'd3,3'd3,3'd2,3'd2,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_28_21[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd2,3'd3,3'd3},
'{3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd1,3'd0,3'd1,3'd0,3'd0},
'{3'd1,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd2,3'd2,3'd1,3'd0,3'd0,3'd1,3'd1}};

parameter bit [2:0] SpriteTableG_28_22[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd4,3'd1,3'd3,3'd3,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd3,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_28_23[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1}};

parameter bit [2:0] SpriteTableG_28_24[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_28_25[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd3,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd3,3'd1,3'd1},
'{3'd0,3'd0,3'd4,3'd1,3'd3,3'd2,3'd1,3'd1},
'{3'd1,3'd3,3'd3,3'd2,3'd1,3'd1,3'd1,3'd1},
'{3'd3,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1}};

parameter bit [2:0] SpriteTableG_28_26[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd2},
'{3'd1,3'd1,3'd1,3'd0,3'd4,3'd0,3'd4,3'd2},
'{3'd1,3'd1,3'd0,3'd4,3'd4,3'd0,3'd1,3'd3},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd2,3'd3},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd4,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd2,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_28_27[7:0][7:0] = '{'{3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd4,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_28_28[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_28_29[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd4,3'd1,3'd4,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd4,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd1,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_28_30[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd2},
'{3'd0,3'd0,3'd0,3'd4,3'd1,3'd0,3'd1,3'd3},
'{3'd0,3'd0,3'd4,3'd1,3'd4,3'd4,3'd4,3'd1},
'{3'd0,3'd0,3'd0,3'd4,3'd4,3'd4,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_28_31[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd2,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd2,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd1,3'd4,3'd0,3'd1,3'd3},
'{3'd0,3'd0,3'd0,3'd1,3'd4,3'd0,3'd0,3'd2},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_28_32[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd4,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_28_33[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_28_34[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0},
'{3'd3,3'd2,3'd2,3'd3,3'd2,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_28_35[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_29_0[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_29_1[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd4,3'd4,3'd4},
'{3'd0,3'd0,3'd4,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd4,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_29_2[7:0][7:0] = '{'{3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd4,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd4,3'd0,3'd0},
'{3'd0,3'd4,3'd4,3'd0,3'd4,3'd1,3'd0,3'd0},
'{3'd4,3'd1,3'd0,3'd0,3'd0,3'd4,3'd0,3'd0},
'{3'd1,3'd4,3'd0,3'd0,3'd0,3'd4,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_29_3[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd4,3'd4,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd0,3'd4,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_29_4[7:0][7:0] = '{'{3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd4,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd1,3'd3,3'd1,3'd4,3'd4,3'd1,3'd3},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd0,3'd0,3'd0,3'd4,3'd1,3'd1,3'd4,3'd0}};

parameter bit [2:0] SpriteTableG_29_5[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_29_6[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0},
'{3'd3,3'd2,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0},
'{3'd3,3'd3,3'd2,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd3,3'd3,3'd3,3'd2,3'd2,3'd2,3'd2,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd2,3'd1,3'd1},
'{3'd3,3'd3,3'd3,3'd2,3'd3,3'd3,3'd1,3'd1}};

parameter bit [2:0] SpriteTableG_29_7[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd0},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1},
'{3'd2,3'd3,3'd3,3'd2,3'd1,3'd2,3'd2,3'd2},
'{3'd1,3'd3,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd3,3'd0,3'd0,3'd0,3'd0,3'd2,3'd3},
'{3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd4,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4}};

parameter bit [2:0] SpriteTableG_29_8[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd4,3'd1,3'd0,3'd3,3'd3,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd3,3'd3,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_29_9[7:0][7:0] = '{'{3'd1,3'd1,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd1},
'{3'd3,3'd3,3'd2,3'd3,3'd2,3'd2,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_29_10[7:0][7:0] = '{'{3'd2,3'd2,3'd1,3'd0,3'd0,3'd1,3'd2,3'd2},
'{3'd0,3'd0,3'd1,3'd2,3'd3,3'd3,3'd3,3'd1},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd2,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd2,3'd0,3'd0,3'd1,3'd0},
'{3'd3,3'd3,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd1,3'd0,3'd1,3'd2,3'd3,3'd2,3'd0},
'{3'd2,3'd2,3'd3,3'd3,3'd3,3'd2,3'd0,3'd1}};

parameter bit [2:0] SpriteTableG_29_11[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd1},
'{3'd3,3'd3,3'd1,3'd0,3'd1,3'd0,3'd1,3'd0},
'{3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd0,3'd0,3'd1,3'd0,3'd0,3'd1,3'd2,3'd2},
'{3'd1,3'd1,3'd0,3'd0,3'd1,3'd1,3'd2,3'd2},
'{3'd1,3'd1,3'd0,3'd1,3'd2,3'd2,3'd2,3'd3},
'{3'd0,3'd0,3'd0,3'd1,3'd2,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_29_12[7:0][7:0] = '{'{3'd0,3'd0,3'd1,3'd2,3'd3,3'd3,3'd2,3'd3},
'{3'd0,3'd1,3'd4,3'd3,3'd3,3'd3,3'd2,3'd3},
'{3'd1,3'd0,3'd4,3'd1,3'd4,3'd1,3'd3,3'd2},
'{3'd1,3'd4,3'd0,3'd0,3'd0,3'd0,3'd2,3'd1},
'{3'd3,3'd3,3'd4,3'd0,3'd4,3'd3,3'd1,3'd0},
'{3'd1,3'd3,3'd4,3'd0,3'd4,3'd3,3'd4,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_29_13[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd4,3'd0,3'd4,3'd3,3'd4,3'd1},
'{3'd3,3'd3,3'd4,3'd0,3'd1,3'd3,3'd2,3'd1},
'{3'd4,3'd4,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1},
'{3'd1,3'd3,3'd0,3'd0,3'd4,3'd1,3'd1,3'd1},
'{3'd1,3'd3,3'd4,3'd0,3'd4,3'd3,3'd1,3'd0}};

parameter bit [2:0] SpriteTableG_29_14[7:0][7:0] = '{'{3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd4,3'd0},
'{3'd1,3'd3,3'd4,3'd0,3'd4,3'd3,3'd2,3'd1},
'{3'd4,3'd1,3'd0,3'd0,3'd0,3'd4,3'd4,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2}};

parameter bit [2:0] SpriteTableG_29_15[7:0][7:0] = '{'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd4,3'd0,3'd2},
'{3'd3,3'd3,3'd4,3'd0,3'd4,3'd3,3'd1,3'd3},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd2,3'd3,3'd3},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd2,3'd3},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd0,3'd0,3'd1,3'd0,3'd0,3'd3,3'd4,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_29_16[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd3,3'd2,3'd2,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd2,3'd2,3'd0,3'd0,3'd0},
'{3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_29_17[7:0][7:0] = '{'{3'd3,3'd2,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd1,3'd0,3'd0},
'{3'd3,3'd2,3'd2,3'd0,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd4,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd3,3'd1,3'd2,3'd1,3'd0,3'd0,3'd1},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd4}};

parameter bit [2:0] SpriteTableG_29_18[7:0][7:0] = '{'{3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_29_19[7:0][7:0] = '{'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1}};

parameter bit [2:0] SpriteTableG_29_20[7:0][7:0] = '{'{3'd2,3'd2,3'd2,3'd1,3'd1,3'd2,3'd2,3'd1},
'{3'd1,3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd0},
'{3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0},
'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0},
'{3'd1,3'd0,3'd1,3'd1,3'd2,3'd2,3'd2,3'd0},
'{3'd1,3'd1,3'd2,3'd2,3'd2,3'd2,3'd2,3'd2},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd3},
'{3'd2,3'd2,3'd2,3'd2,3'd2,3'd1,3'd1,3'd2}};

parameter bit [2:0] SpriteTableG_29_21[7:0][7:0] = '{'{3'd3,3'd2,3'd1,3'd2,3'd3,3'd1,3'd3,3'd3},
'{3'd3,3'd1,3'd2,3'd3,3'd2,3'd1,3'd3,3'd3},
'{3'd3,3'd2,3'd2,3'd3,3'd3,3'd1,3'd4,3'd1},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd0,3'd1},
'{3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd1,3'd3,3'd3,3'd2,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd2,3'd1},
'{3'd1,3'd0,3'd0,3'd1,3'd0,3'd0,3'd1,3'd1}};

parameter bit [2:0] SpriteTableG_29_22[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd1},
'{3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1},
'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd3,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0},
'{3'd4,3'd3,3'd1,3'd0,3'd0,3'd0,3'd2,3'd1}};

parameter bit [2:0] SpriteTableG_29_23[7:0][7:0] = '{'{3'd0,3'd3,3'd2,3'd4,3'd0,3'd1,3'd2,3'd1},
'{3'd0,3'd3,3'd3,3'd3,3'd2,3'd1,3'd1,3'd1},
'{3'd0,3'd3,3'd3,3'd2,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd3,3'd3,3'd2,3'd1,3'd1,3'd1,3'd1},
'{3'd4,3'd3,3'd3,3'd1,3'd0,3'd1,3'd1,3'd1},
'{3'd1,3'd1,3'd2,3'd1,3'd0,3'd1,3'd1,3'd1},
'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_29_24[7:0][7:0] = '{'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd4,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd3,3'd3,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd1,3'd3,3'd3,3'd1,3'd0},
'{3'd1,3'd1,3'd0,3'd2,3'd3,3'd3,3'd3,3'd1},
'{3'd1,3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_29_25[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd0,3'd3,3'd3,3'd3,3'd2,3'd3,3'd3},
'{3'd1,3'd1,3'd3,3'd3,3'd1,3'd0,3'd0,3'd2},
'{3'd1,3'd3,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd3,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_29_26[7:0][7:0] = '{'{3'd2,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd3,3'd3,3'd2,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd1}};

parameter bit [2:0] SpriteTableG_29_27[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_29_28[7:0][7:0] = '{'{3'd3,3'd3,3'd2,3'd2,3'd2,3'd3,3'd3,3'd3},
'{3'd3,3'd2,3'd2,3'd2,3'd2,3'd2,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_29_29[7:0][7:0] = '{'{3'd0,3'd1,3'd1,3'd1,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd1,3'd1,3'd0,3'd4,3'd2,3'd3,3'd3},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd3},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_29_30[7:0][7:0] = '{'{3'd2,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_29_31[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd2,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd2,3'd2,3'd4,3'd0,3'd0,3'd0},
'{3'd3,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_29_32[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_29_33[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_29_34[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_29_35[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_30_0[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_30_1[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd3,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd0,3'd4,3'd1,3'd1,3'd4},
'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_30_2[7:0][7:0] = '{'{3'd0,3'd0,3'd1,3'd4,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4}};

parameter bit [2:0] SpriteTableG_30_3[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd4,3'd4,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd4,3'd3,3'd4},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0},
'{3'd1,3'd0,3'd0,3'd4,3'd1,3'd1,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_30_4[7:0][7:0] = '{'{3'd1,3'd4,3'd1,3'd3,3'd2,3'd0,3'd0,3'd0},
'{3'd1,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd0,3'd0,3'd0},
'{3'd3,3'd2,3'd1,3'd4,3'd1,3'd4,3'd0,3'd0},
'{3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_30_5[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_30_6[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_30_7[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd3,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd3,3'd3,3'd1,3'd1,3'd4,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_30_8[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd4,3'd0},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd0,3'd0,3'd0},
'{3'd2,3'd3,3'd3,3'd3,3'd2,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd1,3'd2,3'd3,3'd0,3'd0,3'd0},
'{3'd4,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_30_9[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0}};

parameter bit [2:0] SpriteTableG_30_10[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd0,3'd0,3'd1,3'd0,3'd0,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd0,3'd1,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_30_11[7:0][7:0] = '{'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd2},
'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd2,3'd3,3'd2},
'{3'd2,3'd2,3'd2,3'd1,3'd2,3'd3,3'd3,3'd2},
'{3'd1,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd1,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3}};

parameter bit [2:0] SpriteTableG_30_12[7:0][7:0] = '{'{3'd3,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd0,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd1,3'd2,3'd2,3'd0,3'd1,3'd3,3'd3,3'd2},
'{3'd0,3'd4,3'd1,3'd0,3'd0,3'd1,3'd3,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_30_13[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd4,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd4},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd2},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd4,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd1,3'd1}};

parameter bit [2:0] SpriteTableG_30_14[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd4,3'd1,3'd0,3'd0,3'd1,3'd4,3'd0},
'{3'd2,3'd4,3'd0,3'd4,3'd2,3'd3,3'd4,3'd0},
'{3'd3,3'd3,3'd2,3'd3,3'd3,3'd3,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_30_15[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd2},
'{3'd2,3'd3,3'd3,3'd3,3'd2,3'd0,3'd0,3'd0},
'{3'd1,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0},
'{3'd1,3'd2,3'd2,3'd2,3'd1,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_30_16[7:0][7:0] = '{'{3'd1,3'd1,3'd2,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0},
'{3'd1,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1},
'{3'd1,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0}};

parameter bit [2:0] SpriteTableG_30_17[7:0][7:0] = '{'{3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd2,3'd1,3'd0,3'd4,3'd2,3'd4,3'd0},
'{3'd0,3'd2,3'd3,3'd2,3'd2,3'd2,3'd0,3'd0},
'{3'd0,3'd2,3'd3,3'd3,3'd3,3'd2,3'd0,3'd0},
'{3'd4,3'd3,3'd3,3'd2,3'd3,3'd2,3'd0,3'd0},
'{3'd2,3'd3,3'd1,3'd0,3'd2,3'd3,3'd1,3'd0},
'{3'd1,3'd2,3'd1,3'd0,3'd1,3'd3,3'd2,3'd4}};

parameter bit [2:0] SpriteTableG_30_18[7:0][7:0] = '{'{3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0}};

parameter bit [2:0] SpriteTableG_30_19[7:0][7:0] = '{'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0},
'{3'd4,3'd0,3'd4,3'd2,3'd2,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd1,3'd2,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd4,3'd2,3'd1,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd1,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_30_20[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd2,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd3,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd2,3'd4,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_30_21[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd3,3'd2,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd2,3'd4,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_30_22[7:0][7:0] = '{'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd1,3'd1,3'd0,3'd1,3'd1,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_30_23[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_30_24[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_30_25[7:0][7:0] = '{'{3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_30_26[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_30_27[7:0][7:0] = '{'{3'd3,3'd3,3'd2,3'd2,3'd1,3'd1,3'd4,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_30_28[7:0][7:0] = '{'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_30_29[7:0][7:0] = '{'{3'd3,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd2,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd3,3'd3,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd4,3'd2,3'd4,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_30_30[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_30_31[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_30_32[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_30_33[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_30_34[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_30_35[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_31_0[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_31_1[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd4,3'd3,3'd4,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_31_2[7:0][7:0] = '{'{3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd3,3'd4,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd3,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd3,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_31_3[7:0][7:0] = '{'{3'd0,3'd4,3'd3,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_31_4[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_31_5[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_31_6[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_31_7[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_31_8[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_31_9[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd1,3'd1},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0},
'{3'd0,3'd1,3'd1,3'd0,3'd0,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_31_10[7:0][7:0] = '{'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_31_11[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd3,3'd3,3'd1,3'd0,3'd1,3'd1,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_31_12[7:0][7:0] = '{'{3'd3,3'd3,3'd3,3'd2,3'd3,3'd2,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0,3'd0},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd4,3'd0,3'd0},
'{3'd3,3'd3,3'd3,3'd3,3'd3,3'd2,3'd0,3'd0},
'{3'd2,3'd3,3'd3,3'd3,3'd3,3'd3,3'd1,3'd0},
'{3'd0,3'd1,3'd3,3'd2,3'd4,3'd4,3'd0,3'd0},
'{3'd0,3'd4,3'd3,3'd4,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_31_13[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd2,3'd2,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_31_14[7:0][7:0] = '{'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_31_15[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_31_16[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0},
'{3'd0,3'd0,3'd1,3'd1,3'd1,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_31_17[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_31_18[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_31_19[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_31_20[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_31_21[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_31_22[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_31_23[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_31_24[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_31_25[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_31_26[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_31_27[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd1,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_31_28[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_31_29[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_31_30[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_31_31[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_31_32[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_31_33[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd4,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_31_34[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

parameter bit [2:0] SpriteTableG_31_35[7:0][7:0] = '{'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0},
'{3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0,3'd0}};

logic [9:0] SpriteTableB;

parameter bit [7:0] SpritePaletteB[3:0] = '{8'd255, 8'd174, 8'd81, 8'd0};

	always_comb
	begin
		SpriteTableB = 10'd0;
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableB = SpriteTableB_0_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableB = SpriteTableB_0_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableB = SpriteTableB_0_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableB = SpriteTableB_0_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableB = SpriteTableB_0_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableB = SpriteTableB_0_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableB = SpriteTableB_0_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableB = SpriteTableB_0_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableB = SpriteTableB_0_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableB = SpriteTableB_0_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableB = SpriteTableB_0_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableB = SpriteTableB_0_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableB = SpriteTableB_0_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_0_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableB = SpriteTableB_0_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableB = SpriteTableB_0_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableB = SpriteTableB_0_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableB = SpriteTableB_0_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableB = SpriteTableB_0_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableB = SpriteTableB_0_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableB = SpriteTableB_0_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableB = SpriteTableB_0_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableB = SpriteTableB_0_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableB = SpriteTableB_0_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableB = SpriteTableB_0_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableB = SpriteTableB_0_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableB = SpriteTableB_0_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableB = SpriteTableB_0_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableB = SpriteTableB_0_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableB = SpriteTableB_0_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableB = SpriteTableB_0_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableB = SpriteTableB_0_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableB = SpriteTableB_0_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableB = SpriteTableB_0_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableB = SpriteTableB_0_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd0 && SpriteX < 10'd8 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableB = SpriteTableB_0_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableB = SpriteTableB_1_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableB = SpriteTableB_1_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableB = SpriteTableB_1_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableB = SpriteTableB_1_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableB = SpriteTableB_1_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableB = SpriteTableB_1_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableB = SpriteTableB_1_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableB = SpriteTableB_1_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableB = SpriteTableB_1_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableB = SpriteTableB_1_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableB = SpriteTableB_1_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableB = SpriteTableB_1_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableB = SpriteTableB_1_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_1_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableB = SpriteTableB_1_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableB = SpriteTableB_1_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableB = SpriteTableB_1_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableB = SpriteTableB_1_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableB = SpriteTableB_1_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableB = SpriteTableB_1_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableB = SpriteTableB_1_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableB = SpriteTableB_1_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableB = SpriteTableB_1_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableB = SpriteTableB_1_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableB = SpriteTableB_1_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableB = SpriteTableB_1_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableB = SpriteTableB_1_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableB = SpriteTableB_1_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableB = SpriteTableB_1_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableB = SpriteTableB_1_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableB = SpriteTableB_1_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableB = SpriteTableB_1_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableB = SpriteTableB_1_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableB = SpriteTableB_1_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableB = SpriteTableB_1_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd8 && SpriteX < 10'd16 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableB = SpriteTableB_1_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableB = SpriteTableB_2_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableB = SpriteTableB_2_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableB = SpriteTableB_2_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableB = SpriteTableB_2_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableB = SpriteTableB_2_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableB = SpriteTableB_2_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableB = SpriteTableB_2_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableB = SpriteTableB_2_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableB = SpriteTableB_2_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableB = SpriteTableB_2_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableB = SpriteTableB_2_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableB = SpriteTableB_2_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableB = SpriteTableB_2_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_2_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableB = SpriteTableB_2_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableB = SpriteTableB_2_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableB = SpriteTableB_2_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableB = SpriteTableB_2_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableB = SpriteTableB_2_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableB = SpriteTableB_2_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableB = SpriteTableB_2_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableB = SpriteTableB_2_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableB = SpriteTableB_2_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableB = SpriteTableB_2_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableB = SpriteTableB_2_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableB = SpriteTableB_2_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableB = SpriteTableB_2_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableB = SpriteTableB_2_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableB = SpriteTableB_2_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableB = SpriteTableB_2_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableB = SpriteTableB_2_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableB = SpriteTableB_2_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableB = SpriteTableB_2_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableB = SpriteTableB_2_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableB = SpriteTableB_2_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd16 && SpriteX < 10'd24 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableB = SpriteTableB_2_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableB = SpriteTableB_3_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableB = SpriteTableB_3_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableB = SpriteTableB_3_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableB = SpriteTableB_3_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableB = SpriteTableB_3_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableB = SpriteTableB_3_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableB = SpriteTableB_3_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableB = SpriteTableB_3_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableB = SpriteTableB_3_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableB = SpriteTableB_3_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableB = SpriteTableB_3_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableB = SpriteTableB_3_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableB = SpriteTableB_3_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_3_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableB = SpriteTableB_3_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableB = SpriteTableB_3_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableB = SpriteTableB_3_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableB = SpriteTableB_3_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableB = SpriteTableB_3_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableB = SpriteTableB_3_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableB = SpriteTableB_3_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableB = SpriteTableB_3_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableB = SpriteTableB_3_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableB = SpriteTableB_3_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableB = SpriteTableB_3_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableB = SpriteTableB_3_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableB = SpriteTableB_3_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableB = SpriteTableB_3_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableB = SpriteTableB_3_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableB = SpriteTableB_3_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableB = SpriteTableB_3_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableB = SpriteTableB_3_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableB = SpriteTableB_3_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableB = SpriteTableB_3_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableB = SpriteTableB_3_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd24 && SpriteX < 10'd32 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableB = SpriteTableB_3_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableB = SpriteTableB_4_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableB = SpriteTableB_4_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableB = SpriteTableB_4_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableB = SpriteTableB_4_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableB = SpriteTableB_4_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableB = SpriteTableB_4_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableB = SpriteTableB_4_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableB = SpriteTableB_4_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableB = SpriteTableB_4_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableB = SpriteTableB_4_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableB = SpriteTableB_4_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableB = SpriteTableB_4_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableB = SpriteTableB_4_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_4_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableB = SpriteTableB_4_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableB = SpriteTableB_4_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableB = SpriteTableB_4_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableB = SpriteTableB_4_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableB = SpriteTableB_4_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableB = SpriteTableB_4_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableB = SpriteTableB_4_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableB = SpriteTableB_4_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableB = SpriteTableB_4_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableB = SpriteTableB_4_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableB = SpriteTableB_4_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableB = SpriteTableB_4_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableB = SpriteTableB_4_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableB = SpriteTableB_4_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableB = SpriteTableB_4_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableB = SpriteTableB_4_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableB = SpriteTableB_4_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableB = SpriteTableB_4_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableB = SpriteTableB_4_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableB = SpriteTableB_4_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableB = SpriteTableB_4_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd32 && SpriteX < 10'd40 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableB = SpriteTableB_4_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableB = SpriteTableB_5_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableB = SpriteTableB_5_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableB = SpriteTableB_5_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableB = SpriteTableB_5_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableB = SpriteTableB_5_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableB = SpriteTableB_5_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableB = SpriteTableB_5_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableB = SpriteTableB_5_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableB = SpriteTableB_5_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableB = SpriteTableB_5_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableB = SpriteTableB_5_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableB = SpriteTableB_5_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableB = SpriteTableB_5_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_5_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableB = SpriteTableB_5_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableB = SpriteTableB_5_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableB = SpriteTableB_5_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableB = SpriteTableB_5_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableB = SpriteTableB_5_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableB = SpriteTableB_5_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableB = SpriteTableB_5_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableB = SpriteTableB_5_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableB = SpriteTableB_5_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableB = SpriteTableB_5_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableB = SpriteTableB_5_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableB = SpriteTableB_5_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableB = SpriteTableB_5_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableB = SpriteTableB_5_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableB = SpriteTableB_5_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableB = SpriteTableB_5_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableB = SpriteTableB_5_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableB = SpriteTableB_5_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableB = SpriteTableB_5_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableB = SpriteTableB_5_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableB = SpriteTableB_5_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd40 && SpriteX < 10'd48 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableB = SpriteTableB_5_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableB = SpriteTableB_6_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableB = SpriteTableB_6_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableB = SpriteTableB_6_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableB = SpriteTableB_6_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableB = SpriteTableB_6_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableB = SpriteTableB_6_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableB = SpriteTableB_6_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableB = SpriteTableB_6_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableB = SpriteTableB_6_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableB = SpriteTableB_6_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableB = SpriteTableB_6_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableB = SpriteTableB_6_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableB = SpriteTableB_6_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_6_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableB = SpriteTableB_6_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableB = SpriteTableB_6_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableB = SpriteTableB_6_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableB = SpriteTableB_6_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableB = SpriteTableB_6_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableB = SpriteTableB_6_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableB = SpriteTableB_6_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableB = SpriteTableB_6_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableB = SpriteTableB_6_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableB = SpriteTableB_6_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableB = SpriteTableB_6_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableB = SpriteTableB_6_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableB = SpriteTableB_6_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableB = SpriteTableB_6_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableB = SpriteTableB_6_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableB = SpriteTableB_6_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableB = SpriteTableB_6_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableB = SpriteTableB_6_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableB = SpriteTableB_6_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableB = SpriteTableB_6_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableB = SpriteTableB_6_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd48 && SpriteX < 10'd56 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableB = SpriteTableB_6_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableB = SpriteTableB_7_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableB = SpriteTableB_7_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableB = SpriteTableB_7_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableB = SpriteTableB_7_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableB = SpriteTableB_7_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableB = SpriteTableB_7_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableB = SpriteTableB_7_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableB = SpriteTableB_7_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableB = SpriteTableB_7_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableB = SpriteTableB_7_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableB = SpriteTableB_7_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableB = SpriteTableB_7_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableB = SpriteTableB_7_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_7_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableB = SpriteTableB_7_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableB = SpriteTableB_7_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableB = SpriteTableB_7_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableB = SpriteTableB_7_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableB = SpriteTableB_7_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableB = SpriteTableB_7_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableB = SpriteTableB_7_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableB = SpriteTableB_7_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableB = SpriteTableB_7_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableB = SpriteTableB_7_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableB = SpriteTableB_7_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableB = SpriteTableB_7_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableB = SpriteTableB_7_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableB = SpriteTableB_7_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableB = SpriteTableB_7_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableB = SpriteTableB_7_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableB = SpriteTableB_7_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableB = SpriteTableB_7_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableB = SpriteTableB_7_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableB = SpriteTableB_7_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableB = SpriteTableB_7_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd56 && SpriteX < 10'd64 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableB = SpriteTableB_7_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableB = SpriteTableB_8_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableB = SpriteTableB_8_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableB = SpriteTableB_8_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableB = SpriteTableB_8_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableB = SpriteTableB_8_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableB = SpriteTableB_8_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableB = SpriteTableB_8_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableB = SpriteTableB_8_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableB = SpriteTableB_8_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableB = SpriteTableB_8_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableB = SpriteTableB_8_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableB = SpriteTableB_8_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableB = SpriteTableB_8_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_8_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableB = SpriteTableB_8_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableB = SpriteTableB_8_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableB = SpriteTableB_8_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableB = SpriteTableB_8_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableB = SpriteTableB_8_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableB = SpriteTableB_8_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableB = SpriteTableB_8_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableB = SpriteTableB_8_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableB = SpriteTableB_8_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableB = SpriteTableB_8_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableB = SpriteTableB_8_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableB = SpriteTableB_8_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableB = SpriteTableB_8_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableB = SpriteTableB_8_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableB = SpriteTableB_8_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableB = SpriteTableB_8_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableB = SpriteTableB_8_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableB = SpriteTableB_8_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableB = SpriteTableB_8_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableB = SpriteTableB_8_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableB = SpriteTableB_8_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd64 && SpriteX < 10'd72 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableB = SpriteTableB_8_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableB = SpriteTableB_9_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableB = SpriteTableB_9_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableB = SpriteTableB_9_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableB = SpriteTableB_9_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableB = SpriteTableB_9_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableB = SpriteTableB_9_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableB = SpriteTableB_9_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableB = SpriteTableB_9_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableB = SpriteTableB_9_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableB = SpriteTableB_9_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableB = SpriteTableB_9_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableB = SpriteTableB_9_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableB = SpriteTableB_9_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_9_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableB = SpriteTableB_9_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableB = SpriteTableB_9_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableB = SpriteTableB_9_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableB = SpriteTableB_9_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableB = SpriteTableB_9_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableB = SpriteTableB_9_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableB = SpriteTableB_9_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableB = SpriteTableB_9_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableB = SpriteTableB_9_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableB = SpriteTableB_9_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableB = SpriteTableB_9_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableB = SpriteTableB_9_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableB = SpriteTableB_9_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableB = SpriteTableB_9_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableB = SpriteTableB_9_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableB = SpriteTableB_9_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableB = SpriteTableB_9_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableB = SpriteTableB_9_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableB = SpriteTableB_9_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableB = SpriteTableB_9_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableB = SpriteTableB_9_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd72 && SpriteX < 10'd80 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableB = SpriteTableB_9_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableB = SpriteTableB_10_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableB = SpriteTableB_10_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableB = SpriteTableB_10_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableB = SpriteTableB_10_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableB = SpriteTableB_10_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableB = SpriteTableB_10_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableB = SpriteTableB_10_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableB = SpriteTableB_10_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableB = SpriteTableB_10_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableB = SpriteTableB_10_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableB = SpriteTableB_10_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableB = SpriteTableB_10_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableB = SpriteTableB_10_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_10_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableB = SpriteTableB_10_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableB = SpriteTableB_10_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableB = SpriteTableB_10_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableB = SpriteTableB_10_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableB = SpriteTableB_10_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableB = SpriteTableB_10_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableB = SpriteTableB_10_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableB = SpriteTableB_10_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableB = SpriteTableB_10_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableB = SpriteTableB_10_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableB = SpriteTableB_10_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableB = SpriteTableB_10_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableB = SpriteTableB_10_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableB = SpriteTableB_10_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableB = SpriteTableB_10_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableB = SpriteTableB_10_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableB = SpriteTableB_10_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableB = SpriteTableB_10_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableB = SpriteTableB_10_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableB = SpriteTableB_10_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableB = SpriteTableB_10_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd80 && SpriteX < 10'd88 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableB = SpriteTableB_10_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableB = SpriteTableB_11_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableB = SpriteTableB_11_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableB = SpriteTableB_11_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableB = SpriteTableB_11_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableB = SpriteTableB_11_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableB = SpriteTableB_11_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableB = SpriteTableB_11_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableB = SpriteTableB_11_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableB = SpriteTableB_11_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableB = SpriteTableB_11_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableB = SpriteTableB_11_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableB = SpriteTableB_11_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableB = SpriteTableB_11_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_11_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableB = SpriteTableB_11_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableB = SpriteTableB_11_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableB = SpriteTableB_11_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableB = SpriteTableB_11_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableB = SpriteTableB_11_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableB = SpriteTableB_11_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableB = SpriteTableB_11_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableB = SpriteTableB_11_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableB = SpriteTableB_11_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableB = SpriteTableB_11_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableB = SpriteTableB_11_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableB = SpriteTableB_11_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableB = SpriteTableB_11_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableB = SpriteTableB_11_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableB = SpriteTableB_11_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableB = SpriteTableB_11_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableB = SpriteTableB_11_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableB = SpriteTableB_11_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableB = SpriteTableB_11_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableB = SpriteTableB_11_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableB = SpriteTableB_11_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd88 && SpriteX < 10'd96 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableB = SpriteTableB_11_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableB = SpriteTableB_12_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableB = SpriteTableB_12_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableB = SpriteTableB_12_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableB = SpriteTableB_12_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableB = SpriteTableB_12_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableB = SpriteTableB_12_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableB = SpriteTableB_12_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableB = SpriteTableB_12_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableB = SpriteTableB_12_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableB = SpriteTableB_12_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableB = SpriteTableB_12_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableB = SpriteTableB_12_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableB = SpriteTableB_12_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_12_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableB = SpriteTableB_12_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableB = SpriteTableB_12_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableB = SpriteTableB_12_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableB = SpriteTableB_12_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableB = SpriteTableB_12_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableB = SpriteTableB_12_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableB = SpriteTableB_12_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableB = SpriteTableB_12_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableB = SpriteTableB_12_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableB = SpriteTableB_12_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableB = SpriteTableB_12_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableB = SpriteTableB_12_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableB = SpriteTableB_12_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableB = SpriteTableB_12_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableB = SpriteTableB_12_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableB = SpriteTableB_12_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableB = SpriteTableB_12_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableB = SpriteTableB_12_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableB = SpriteTableB_12_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableB = SpriteTableB_12_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableB = SpriteTableB_12_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd96 && SpriteX < 10'd104 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableB = SpriteTableB_12_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableB = SpriteTableB_13_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableB = SpriteTableB_13_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableB = SpriteTableB_13_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableB = SpriteTableB_13_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableB = SpriteTableB_13_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableB = SpriteTableB_13_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableB = SpriteTableB_13_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableB = SpriteTableB_13_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableB = SpriteTableB_13_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableB = SpriteTableB_13_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableB = SpriteTableB_13_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableB = SpriteTableB_13_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableB = SpriteTableB_13_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_13_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableB = SpriteTableB_13_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableB = SpriteTableB_13_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableB = SpriteTableB_13_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableB = SpriteTableB_13_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableB = SpriteTableB_13_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableB = SpriteTableB_13_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableB = SpriteTableB_13_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableB = SpriteTableB_13_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableB = SpriteTableB_13_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableB = SpriteTableB_13_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableB = SpriteTableB_13_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableB = SpriteTableB_13_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableB = SpriteTableB_13_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableB = SpriteTableB_13_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableB = SpriteTableB_13_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableB = SpriteTableB_13_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableB = SpriteTableB_13_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableB = SpriteTableB_13_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableB = SpriteTableB_13_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableB = SpriteTableB_13_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableB = SpriteTableB_13_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd104 && SpriteX < 10'd112 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableB = SpriteTableB_13_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableB = SpriteTableB_14_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableB = SpriteTableB_14_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableB = SpriteTableB_14_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableB = SpriteTableB_14_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableB = SpriteTableB_14_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableB = SpriteTableB_14_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableB = SpriteTableB_14_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableB = SpriteTableB_14_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableB = SpriteTableB_14_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableB = SpriteTableB_14_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableB = SpriteTableB_14_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableB = SpriteTableB_14_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableB = SpriteTableB_14_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_14_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableB = SpriteTableB_14_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableB = SpriteTableB_14_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableB = SpriteTableB_14_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableB = SpriteTableB_14_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableB = SpriteTableB_14_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableB = SpriteTableB_14_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableB = SpriteTableB_14_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableB = SpriteTableB_14_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableB = SpriteTableB_14_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableB = SpriteTableB_14_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableB = SpriteTableB_14_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableB = SpriteTableB_14_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableB = SpriteTableB_14_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableB = SpriteTableB_14_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableB = SpriteTableB_14_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableB = SpriteTableB_14_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableB = SpriteTableB_14_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableB = SpriteTableB_14_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableB = SpriteTableB_14_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableB = SpriteTableB_14_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableB = SpriteTableB_14_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd112 && SpriteX < 10'd120 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableB = SpriteTableB_14_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableB = SpriteTableB_15_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableB = SpriteTableB_15_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableB = SpriteTableB_15_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableB = SpriteTableB_15_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableB = SpriteTableB_15_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableB = SpriteTableB_15_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableB = SpriteTableB_15_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableB = SpriteTableB_15_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableB = SpriteTableB_15_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableB = SpriteTableB_15_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableB = SpriteTableB_15_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableB = SpriteTableB_15_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableB = SpriteTableB_15_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_15_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableB = SpriteTableB_15_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableB = SpriteTableB_15_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableB = SpriteTableB_15_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableB = SpriteTableB_15_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableB = SpriteTableB_15_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableB = SpriteTableB_15_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableB = SpriteTableB_15_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableB = SpriteTableB_15_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableB = SpriteTableB_15_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableB = SpriteTableB_15_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableB = SpriteTableB_15_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableB = SpriteTableB_15_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableB = SpriteTableB_15_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableB = SpriteTableB_15_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableB = SpriteTableB_15_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableB = SpriteTableB_15_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableB = SpriteTableB_15_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableB = SpriteTableB_15_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableB = SpriteTableB_15_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableB = SpriteTableB_15_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableB = SpriteTableB_15_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd120 && SpriteX < 10'd128 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableB = SpriteTableB_15_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableB = SpriteTableB_16_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableB = SpriteTableB_16_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableB = SpriteTableB_16_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableB = SpriteTableB_16_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableB = SpriteTableB_16_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableB = SpriteTableB_16_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableB = SpriteTableB_16_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableB = SpriteTableB_16_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableB = SpriteTableB_16_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableB = SpriteTableB_16_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableB = SpriteTableB_16_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableB = SpriteTableB_16_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableB = SpriteTableB_16_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_16_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableB = SpriteTableB_16_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableB = SpriteTableB_16_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableB = SpriteTableB_16_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableB = SpriteTableB_16_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableB = SpriteTableB_16_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableB = SpriteTableB_16_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableB = SpriteTableB_16_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableB = SpriteTableB_16_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableB = SpriteTableB_16_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableB = SpriteTableB_16_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableB = SpriteTableB_16_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableB = SpriteTableB_16_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableB = SpriteTableB_16_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableB = SpriteTableB_16_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableB = SpriteTableB_16_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableB = SpriteTableB_16_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableB = SpriteTableB_16_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableB = SpriteTableB_16_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableB = SpriteTableB_16_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableB = SpriteTableB_16_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableB = SpriteTableB_16_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd128 && SpriteX < 10'd136 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableB = SpriteTableB_16_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableB = SpriteTableB_17_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableB = SpriteTableB_17_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableB = SpriteTableB_17_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableB = SpriteTableB_17_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableB = SpriteTableB_17_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableB = SpriteTableB_17_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableB = SpriteTableB_17_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableB = SpriteTableB_17_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableB = SpriteTableB_17_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableB = SpriteTableB_17_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableB = SpriteTableB_17_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableB = SpriteTableB_17_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableB = SpriteTableB_17_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_17_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableB = SpriteTableB_17_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableB = SpriteTableB_17_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableB = SpriteTableB_17_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableB = SpriteTableB_17_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableB = SpriteTableB_17_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableB = SpriteTableB_17_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableB = SpriteTableB_17_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableB = SpriteTableB_17_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableB = SpriteTableB_17_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableB = SpriteTableB_17_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableB = SpriteTableB_17_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableB = SpriteTableB_17_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableB = SpriteTableB_17_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableB = SpriteTableB_17_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableB = SpriteTableB_17_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableB = SpriteTableB_17_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableB = SpriteTableB_17_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableB = SpriteTableB_17_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableB = SpriteTableB_17_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableB = SpriteTableB_17_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableB = SpriteTableB_17_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd136 && SpriteX < 10'd144 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableB = SpriteTableB_17_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableB = SpriteTableB_18_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableB = SpriteTableB_18_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableB = SpriteTableB_18_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableB = SpriteTableB_18_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableB = SpriteTableB_18_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableB = SpriteTableB_18_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableB = SpriteTableB_18_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableB = SpriteTableB_18_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableB = SpriteTableB_18_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableB = SpriteTableB_18_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableB = SpriteTableB_18_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableB = SpriteTableB_18_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableB = SpriteTableB_18_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_18_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableB = SpriteTableB_18_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableB = SpriteTableB_18_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableB = SpriteTableB_18_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableB = SpriteTableB_18_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableB = SpriteTableB_18_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableB = SpriteTableB_18_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableB = SpriteTableB_18_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableB = SpriteTableB_18_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableB = SpriteTableB_18_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableB = SpriteTableB_18_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableB = SpriteTableB_18_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableB = SpriteTableB_18_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableB = SpriteTableB_18_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableB = SpriteTableB_18_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableB = SpriteTableB_18_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableB = SpriteTableB_18_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableB = SpriteTableB_18_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableB = SpriteTableB_18_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableB = SpriteTableB_18_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableB = SpriteTableB_18_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableB = SpriteTableB_18_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd144 && SpriteX < 10'd152 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableB = SpriteTableB_18_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableB = SpriteTableB_19_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableB = SpriteTableB_19_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableB = SpriteTableB_19_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableB = SpriteTableB_19_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableB = SpriteTableB_19_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableB = SpriteTableB_19_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableB = SpriteTableB_19_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableB = SpriteTableB_19_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableB = SpriteTableB_19_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableB = SpriteTableB_19_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableB = SpriteTableB_19_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableB = SpriteTableB_19_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableB = SpriteTableB_19_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_19_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableB = SpriteTableB_19_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableB = SpriteTableB_19_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableB = SpriteTableB_19_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableB = SpriteTableB_19_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableB = SpriteTableB_19_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableB = SpriteTableB_19_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableB = SpriteTableB_19_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableB = SpriteTableB_19_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableB = SpriteTableB_19_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableB = SpriteTableB_19_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableB = SpriteTableB_19_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableB = SpriteTableB_19_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableB = SpriteTableB_19_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableB = SpriteTableB_19_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableB = SpriteTableB_19_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableB = SpriteTableB_19_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableB = SpriteTableB_19_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableB = SpriteTableB_19_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableB = SpriteTableB_19_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableB = SpriteTableB_19_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableB = SpriteTableB_19_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd152 && SpriteX < 10'd160 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableB = SpriteTableB_19_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableB = SpriteTableB_20_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableB = SpriteTableB_20_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableB = SpriteTableB_20_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableB = SpriteTableB_20_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableB = SpriteTableB_20_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableB = SpriteTableB_20_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableB = SpriteTableB_20_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableB = SpriteTableB_20_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableB = SpriteTableB_20_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableB = SpriteTableB_20_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableB = SpriteTableB_20_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableB = SpriteTableB_20_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableB = SpriteTableB_20_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_20_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableB = SpriteTableB_20_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableB = SpriteTableB_20_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableB = SpriteTableB_20_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableB = SpriteTableB_20_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableB = SpriteTableB_20_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableB = SpriteTableB_20_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableB = SpriteTableB_20_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableB = SpriteTableB_20_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableB = SpriteTableB_20_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableB = SpriteTableB_20_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableB = SpriteTableB_20_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableB = SpriteTableB_20_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableB = SpriteTableB_20_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableB = SpriteTableB_20_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableB = SpriteTableB_20_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableB = SpriteTableB_20_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableB = SpriteTableB_20_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableB = SpriteTableB_20_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableB = SpriteTableB_20_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableB = SpriteTableB_20_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableB = SpriteTableB_20_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd160 && SpriteX < 10'd168 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableB = SpriteTableB_20_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableB = SpriteTableB_21_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableB = SpriteTableB_21_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableB = SpriteTableB_21_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableB = SpriteTableB_21_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableB = SpriteTableB_21_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableB = SpriteTableB_21_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableB = SpriteTableB_21_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableB = SpriteTableB_21_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableB = SpriteTableB_21_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableB = SpriteTableB_21_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableB = SpriteTableB_21_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableB = SpriteTableB_21_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableB = SpriteTableB_21_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_21_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableB = SpriteTableB_21_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableB = SpriteTableB_21_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableB = SpriteTableB_21_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableB = SpriteTableB_21_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableB = SpriteTableB_21_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableB = SpriteTableB_21_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableB = SpriteTableB_21_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableB = SpriteTableB_21_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableB = SpriteTableB_21_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableB = SpriteTableB_21_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableB = SpriteTableB_21_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableB = SpriteTableB_21_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableB = SpriteTableB_21_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableB = SpriteTableB_21_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableB = SpriteTableB_21_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableB = SpriteTableB_21_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableB = SpriteTableB_21_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableB = SpriteTableB_21_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableB = SpriteTableB_21_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableB = SpriteTableB_21_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableB = SpriteTableB_21_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd168 && SpriteX < 10'd176 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableB = SpriteTableB_21_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableB = SpriteTableB_22_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableB = SpriteTableB_22_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableB = SpriteTableB_22_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableB = SpriteTableB_22_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableB = SpriteTableB_22_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableB = SpriteTableB_22_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableB = SpriteTableB_22_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableB = SpriteTableB_22_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableB = SpriteTableB_22_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableB = SpriteTableB_22_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableB = SpriteTableB_22_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableB = SpriteTableB_22_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableB = SpriteTableB_22_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_22_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableB = SpriteTableB_22_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableB = SpriteTableB_22_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableB = SpriteTableB_22_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableB = SpriteTableB_22_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableB = SpriteTableB_22_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableB = SpriteTableB_22_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableB = SpriteTableB_22_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableB = SpriteTableB_22_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableB = SpriteTableB_22_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableB = SpriteTableB_22_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableB = SpriteTableB_22_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableB = SpriteTableB_22_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableB = SpriteTableB_22_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableB = SpriteTableB_22_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableB = SpriteTableB_22_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableB = SpriteTableB_22_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableB = SpriteTableB_22_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableB = SpriteTableB_22_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableB = SpriteTableB_22_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableB = SpriteTableB_22_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableB = SpriteTableB_22_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd176 && SpriteX < 10'd184 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableB = SpriteTableB_22_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableB = SpriteTableB_23_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableB = SpriteTableB_23_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableB = SpriteTableB_23_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableB = SpriteTableB_23_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableB = SpriteTableB_23_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableB = SpriteTableB_23_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableB = SpriteTableB_23_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableB = SpriteTableB_23_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableB = SpriteTableB_23_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableB = SpriteTableB_23_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableB = SpriteTableB_23_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableB = SpriteTableB_23_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableB = SpriteTableB_23_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_23_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableB = SpriteTableB_23_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableB = SpriteTableB_23_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableB = SpriteTableB_23_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableB = SpriteTableB_23_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableB = SpriteTableB_23_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableB = SpriteTableB_23_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableB = SpriteTableB_23_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableB = SpriteTableB_23_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableB = SpriteTableB_23_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableB = SpriteTableB_23_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableB = SpriteTableB_23_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableB = SpriteTableB_23_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableB = SpriteTableB_23_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableB = SpriteTableB_23_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableB = SpriteTableB_23_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableB = SpriteTableB_23_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableB = SpriteTableB_23_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableB = SpriteTableB_23_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableB = SpriteTableB_23_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableB = SpriteTableB_23_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableB = SpriteTableB_23_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd184 && SpriteX < 10'd192 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableB = SpriteTableB_23_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableB = SpriteTableB_24_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableB = SpriteTableB_24_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableB = SpriteTableB_24_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableB = SpriteTableB_24_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableB = SpriteTableB_24_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableB = SpriteTableB_24_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableB = SpriteTableB_24_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableB = SpriteTableB_24_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableB = SpriteTableB_24_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableB = SpriteTableB_24_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableB = SpriteTableB_24_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableB = SpriteTableB_24_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableB = SpriteTableB_24_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_24_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableB = SpriteTableB_24_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableB = SpriteTableB_24_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableB = SpriteTableB_24_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableB = SpriteTableB_24_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableB = SpriteTableB_24_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableB = SpriteTableB_24_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableB = SpriteTableB_24_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableB = SpriteTableB_24_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableB = SpriteTableB_24_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableB = SpriteTableB_24_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableB = SpriteTableB_24_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableB = SpriteTableB_24_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableB = SpriteTableB_24_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableB = SpriteTableB_24_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableB = SpriteTableB_24_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableB = SpriteTableB_24_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableB = SpriteTableB_24_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableB = SpriteTableB_24_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableB = SpriteTableB_24_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableB = SpriteTableB_24_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableB = SpriteTableB_24_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd192 && SpriteX < 10'd200 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableB = SpriteTableB_24_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableB = SpriteTableB_25_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableB = SpriteTableB_25_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableB = SpriteTableB_25_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableB = SpriteTableB_25_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableB = SpriteTableB_25_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableB = SpriteTableB_25_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableB = SpriteTableB_25_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableB = SpriteTableB_25_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableB = SpriteTableB_25_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableB = SpriteTableB_25_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableB = SpriteTableB_25_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableB = SpriteTableB_25_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableB = SpriteTableB_25_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_25_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableB = SpriteTableB_25_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableB = SpriteTableB_25_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableB = SpriteTableB_25_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableB = SpriteTableB_25_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableB = SpriteTableB_25_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableB = SpriteTableB_25_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableB = SpriteTableB_25_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableB = SpriteTableB_25_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableB = SpriteTableB_25_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableB = SpriteTableB_25_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableB = SpriteTableB_25_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableB = SpriteTableB_25_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableB = SpriteTableB_25_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableB = SpriteTableB_25_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableB = SpriteTableB_25_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableB = SpriteTableB_25_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableB = SpriteTableB_25_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableB = SpriteTableB_25_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableB = SpriteTableB_25_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableB = SpriteTableB_25_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableB = SpriteTableB_25_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd200 && SpriteX < 10'd208 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableB = SpriteTableB_25_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableB = SpriteTableB_26_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableB = SpriteTableB_26_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableB = SpriteTableB_26_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableB = SpriteTableB_26_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableB = SpriteTableB_26_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableB = SpriteTableB_26_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableB = SpriteTableB_26_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableB = SpriteTableB_26_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableB = SpriteTableB_26_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableB = SpriteTableB_26_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableB = SpriteTableB_26_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableB = SpriteTableB_26_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableB = SpriteTableB_26_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_26_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableB = SpriteTableB_26_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableB = SpriteTableB_26_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableB = SpriteTableB_26_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableB = SpriteTableB_26_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableB = SpriteTableB_26_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableB = SpriteTableB_26_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableB = SpriteTableB_26_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableB = SpriteTableB_26_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableB = SpriteTableB_26_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableB = SpriteTableB_26_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableB = SpriteTableB_26_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableB = SpriteTableB_26_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableB = SpriteTableB_26_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableB = SpriteTableB_26_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableB = SpriteTableB_26_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableB = SpriteTableB_26_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableB = SpriteTableB_26_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableB = SpriteTableB_26_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableB = SpriteTableB_26_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableB = SpriteTableB_26_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableB = SpriteTableB_26_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd208 && SpriteX < 10'd216 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableB = SpriteTableB_26_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableB = SpriteTableB_27_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableB = SpriteTableB_27_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableB = SpriteTableB_27_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableB = SpriteTableB_27_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableB = SpriteTableB_27_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableB = SpriteTableB_27_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableB = SpriteTableB_27_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableB = SpriteTableB_27_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableB = SpriteTableB_27_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableB = SpriteTableB_27_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableB = SpriteTableB_27_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableB = SpriteTableB_27_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableB = SpriteTableB_27_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_27_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableB = SpriteTableB_27_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableB = SpriteTableB_27_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableB = SpriteTableB_27_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableB = SpriteTableB_27_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableB = SpriteTableB_27_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableB = SpriteTableB_27_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableB = SpriteTableB_27_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableB = SpriteTableB_27_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableB = SpriteTableB_27_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableB = SpriteTableB_27_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableB = SpriteTableB_27_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableB = SpriteTableB_27_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableB = SpriteTableB_27_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableB = SpriteTableB_27_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableB = SpriteTableB_27_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableB = SpriteTableB_27_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableB = SpriteTableB_27_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableB = SpriteTableB_27_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableB = SpriteTableB_27_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableB = SpriteTableB_27_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableB = SpriteTableB_27_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd216 && SpriteX < 10'd224 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableB = SpriteTableB_27_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableB = SpriteTableB_28_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableB = SpriteTableB_28_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableB = SpriteTableB_28_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableB = SpriteTableB_28_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableB = SpriteTableB_28_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableB = SpriteTableB_28_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableB = SpriteTableB_28_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableB = SpriteTableB_28_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableB = SpriteTableB_28_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableB = SpriteTableB_28_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableB = SpriteTableB_28_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableB = SpriteTableB_28_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableB = SpriteTableB_28_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_28_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableB = SpriteTableB_28_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableB = SpriteTableB_28_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableB = SpriteTableB_28_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableB = SpriteTableB_28_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableB = SpriteTableB_28_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableB = SpriteTableB_28_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableB = SpriteTableB_28_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableB = SpriteTableB_28_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableB = SpriteTableB_28_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableB = SpriteTableB_28_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableB = SpriteTableB_28_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableB = SpriteTableB_28_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableB = SpriteTableB_28_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableB = SpriteTableB_28_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableB = SpriteTableB_28_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableB = SpriteTableB_28_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableB = SpriteTableB_28_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableB = SpriteTableB_28_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableB = SpriteTableB_28_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableB = SpriteTableB_28_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableB = SpriteTableB_28_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd224 && SpriteX < 10'd232 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableB = SpriteTableB_28_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableB = SpriteTableB_29_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableB = SpriteTableB_29_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableB = SpriteTableB_29_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableB = SpriteTableB_29_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableB = SpriteTableB_29_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableB = SpriteTableB_29_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableB = SpriteTableB_29_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableB = SpriteTableB_29_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableB = SpriteTableB_29_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableB = SpriteTableB_29_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableB = SpriteTableB_29_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableB = SpriteTableB_29_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableB = SpriteTableB_29_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_29_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableB = SpriteTableB_29_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableB = SpriteTableB_29_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableB = SpriteTableB_29_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableB = SpriteTableB_29_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableB = SpriteTableB_29_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableB = SpriteTableB_29_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableB = SpriteTableB_29_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableB = SpriteTableB_29_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableB = SpriteTableB_29_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableB = SpriteTableB_29_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableB = SpriteTableB_29_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableB = SpriteTableB_29_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableB = SpriteTableB_29_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableB = SpriteTableB_29_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableB = SpriteTableB_29_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableB = SpriteTableB_29_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableB = SpriteTableB_29_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableB = SpriteTableB_29_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableB = SpriteTableB_29_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableB = SpriteTableB_29_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableB = SpriteTableB_29_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd232 && SpriteX < 10'd240 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableB = SpriteTableB_29_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableB = SpriteTableB_30_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableB = SpriteTableB_30_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableB = SpriteTableB_30_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableB = SpriteTableB_30_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableB = SpriteTableB_30_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableB = SpriteTableB_30_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableB = SpriteTableB_30_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableB = SpriteTableB_30_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableB = SpriteTableB_30_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableB = SpriteTableB_30_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableB = SpriteTableB_30_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableB = SpriteTableB_30_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableB = SpriteTableB_30_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_30_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableB = SpriteTableB_30_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableB = SpriteTableB_30_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableB = SpriteTableB_30_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableB = SpriteTableB_30_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableB = SpriteTableB_30_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableB = SpriteTableB_30_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableB = SpriteTableB_30_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableB = SpriteTableB_30_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableB = SpriteTableB_30_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableB = SpriteTableB_30_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableB = SpriteTableB_30_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableB = SpriteTableB_30_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableB = SpriteTableB_30_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableB = SpriteTableB_30_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableB = SpriteTableB_30_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableB = SpriteTableB_30_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableB = SpriteTableB_30_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableB = SpriteTableB_30_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableB = SpriteTableB_30_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableB = SpriteTableB_30_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableB = SpriteTableB_30_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd240 && SpriteX < 10'd248 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableB = SpriteTableB_30_35[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd0 && SpriteY < 10'd8)
		begin
		    SpriteTableB = SpriteTableB_31_0[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd8 && SpriteY < 10'd16)
		begin
		    SpriteTableB = SpriteTableB_31_1[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd16 && SpriteY < 10'd24)
		begin
		    SpriteTableB = SpriteTableB_31_2[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd24 && SpriteY < 10'd32)
		begin
		    SpriteTableB = SpriteTableB_31_3[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd32 && SpriteY < 10'd40)
		begin
		    SpriteTableB = SpriteTableB_31_4[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd40 && SpriteY < 10'd48)
		begin
		    SpriteTableB = SpriteTableB_31_5[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd48 && SpriteY < 10'd56)
		begin
		    SpriteTableB = SpriteTableB_31_6[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd56 && SpriteY < 10'd64)
		begin
		    SpriteTableB = SpriteTableB_31_7[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd64 && SpriteY < 10'd72)
		begin
		    SpriteTableB = SpriteTableB_31_8[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd72 && SpriteY < 10'd80)
		begin
		    SpriteTableB = SpriteTableB_31_9[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd80 && SpriteY < 10'd88)
		begin
		    SpriteTableB = SpriteTableB_31_10[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd88 && SpriteY < 10'd96)
		begin
		    SpriteTableB = SpriteTableB_31_11[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd96 && SpriteY < 10'd104)
		begin
		    SpriteTableB = SpriteTableB_31_12[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd104 && SpriteY < 10'd112)
		begin
		    SpriteTableB = SpriteTableB_31_13[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd112 && SpriteY < 10'd120)
		begin
		    SpriteTableB = SpriteTableB_31_14[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd120 && SpriteY < 10'd128)
		begin
		    SpriteTableB = SpriteTableB_31_15[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd128 && SpriteY < 10'd136)
		begin
		    SpriteTableB = SpriteTableB_31_16[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd136 && SpriteY < 10'd144)
		begin
		    SpriteTableB = SpriteTableB_31_17[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd144 && SpriteY < 10'd152)
		begin
		    SpriteTableB = SpriteTableB_31_18[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd152 && SpriteY < 10'd160)
		begin
		    SpriteTableB = SpriteTableB_31_19[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd160 && SpriteY < 10'd168)
		begin
		    SpriteTableB = SpriteTableB_31_20[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd168 && SpriteY < 10'd176)
		begin
		    SpriteTableB = SpriteTableB_31_21[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd176 && SpriteY < 10'd184)
		begin
		    SpriteTableB = SpriteTableB_31_22[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd184 && SpriteY < 10'd192)
		begin
		    SpriteTableB = SpriteTableB_31_23[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd192 && SpriteY < 10'd200)
		begin
		    SpriteTableB = SpriteTableB_31_24[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd200 && SpriteY < 10'd208)
		begin
		    SpriteTableB = SpriteTableB_31_25[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd208 && SpriteY < 10'd216)
		begin
		    SpriteTableB = SpriteTableB_31_26[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd216 && SpriteY < 10'd224)
		begin
		    SpriteTableB = SpriteTableB_31_27[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd224 && SpriteY < 10'd232)
		begin
		    SpriteTableB = SpriteTableB_31_28[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd232 && SpriteY < 10'd240)
		begin
		    SpriteTableB = SpriteTableB_31_29[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd240 && SpriteY < 10'd248)
		begin
		    SpriteTableB = SpriteTableB_31_30[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd248 && SpriteY < 10'd256)
		begin
		    SpriteTableB = SpriteTableB_31_31[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd256 && SpriteY < 10'd264)
		begin
		    SpriteTableB = SpriteTableB_31_32[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd264 && SpriteY < 10'd272)
		begin
		    SpriteTableB = SpriteTableB_31_33[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd272 && SpriteY < 10'd280)
		begin
		    SpriteTableB = SpriteTableB_31_34[Y_Index][X_Index];
		end
		else
		if(SpriteX >= 10'd248 && SpriteX < 10'd256 && SpriteY >= 10'd280 && SpriteY < 10'd288)
		begin
		    SpriteTableB = SpriteTableB_31_35[Y_Index][X_Index];
		end
	end

parameter bit [1:0] SpriteTableB_0_0[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_0_1[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_0_2[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_0_3[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_0_4[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_0_5[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_0_6[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_0_7[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_0_8[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd2}};

parameter bit [1:0] SpriteTableB_0_9[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd1,2'd2,2'd2,2'd2,2'd2}};

parameter bit [1:0] SpriteTableB_0_10[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_0_11[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_0_12[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_0_13[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_0_14[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_0_15[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_0_16[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_0_17[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_0_18[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3}};

parameter bit [1:0] SpriteTableB_0_19[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd1,2'd2,2'd2,2'd2,2'd3},
'{2'd3,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_0_20[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_0_21[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_0_22[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_0_23[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2}};

parameter bit [1:0] SpriteTableB_0_24[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd1,2'd3,2'd2,2'd2,2'd1,2'd1},
'{2'd3,2'd1,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_0_25[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_0_26[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd1,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_0_27[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_0_28[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_0_29[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_0_30[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_0_31[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_0_32[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_0_33[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_0_34[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_0_35[7:0][7:0] = '{'{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1},
'{2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_1_0[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_1_1[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_1_2[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_1_3[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_1_4[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_1_5[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd1},
'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_1_6[7:0][7:0] = '{'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_1_7[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_1_8[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd3,2'd1,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_1_9[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd2,2'd1,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd3,2'd1,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd1,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd1},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2}};

parameter bit [1:0] SpriteTableB_1_10[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd1,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd1,2'd2,2'd2,2'd2,2'd2}};

parameter bit [1:0] SpriteTableB_1_11[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_1_12[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_1_13[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_1_14[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_1_15[7:0][7:0] = '{'{2'd3,2'd3,2'd2,2'd3,2'd2,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_1_16[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_1_17[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd2,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd1},
'{2'd1,2'd2,2'd2,2'd3,2'd3,2'd2,2'd2,2'd2},
'{2'd3,2'd2,2'd2,2'd3,2'd3,2'd2,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_1_18[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd1,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd2,2'd3},
'{2'd3,2'd3,2'd1,2'd2,2'd3,2'd2,2'd2,2'd3},
'{2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_1_19[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd1,2'd2,2'd2,2'd2,2'd2,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd1,2'd3,2'd3,2'd2},
'{2'd1,2'd1,2'd3,2'd3,2'd1,2'd1,2'd3,2'd1},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd2,2'd2,2'd3}};

parameter bit [1:0] SpriteTableB_1_20[7:0][7:0] = '{'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd1,2'd1,2'd3,2'd1,2'd2,2'd3,2'd3},
'{2'd3,2'd1,2'd2,2'd1,2'd2,2'd2,2'd3,2'd1},
'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd1,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_1_21[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_1_22[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_1_23[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd1,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_1_24[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd3},
'{2'd2,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd1},
'{2'd2,2'd3,2'd2,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_1_25[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3}};

parameter bit [1:0] SpriteTableB_1_26[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_1_27[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_1_28[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_1_29[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_1_30[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_1_31[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd2,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_1_32[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd2,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_1_33[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_1_34[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_1_35[7:0][7:0] = '{'{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_2_0[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_2_1[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_2_2[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_2_3[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_2_4[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_2_5[7:0][7:0] = '{'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_2_6[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_2_7[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_2_8[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_2_9[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd2},
'{2'd3,2'd1,2'd1,2'd1,2'd3,2'd3,2'd2,2'd2},
'{2'd2,2'd2,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2}};

parameter bit [1:0] SpriteTableB_2_10[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1},
'{2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_2_11[7:0][7:0] = '{'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_2_12[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd1,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_2_13[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_2_14[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_2_15[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd2,2'd3,2'd2,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd3,2'd2}};

parameter bit [1:0] SpriteTableB_2_16[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_2_17[7:0][7:0] = '{'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd1,2'd3,2'd3,2'd1,2'd3,2'd2,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_2_18[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd2,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd2,2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_2_19[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd2,2'd2,2'd2,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd2,2'd2,2'd2,2'd3},
'{2'd1,2'd3,2'd1,2'd2,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd3,2'd2}};

parameter bit [1:0] SpriteTableB_2_20[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd1},
'{2'd1,2'd3,2'd3,2'd1,2'd3,2'd1,2'd3,2'd2},
'{2'd1,2'd3,2'd3,2'd1,2'd3,2'd1,2'd1,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd2},
'{2'd1,2'd3,2'd3,2'd1,2'd3,2'd2,2'd2,2'd2}};

parameter bit [1:0] SpriteTableB_2_21[7:0][7:0] = '{'{2'd1,2'd3,2'd3,2'd1,2'd3,2'd2,2'd2,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd1,2'd3,2'd1,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3}};

parameter bit [1:0] SpriteTableB_2_22[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd2},
'{2'd1,2'd3,2'd3,2'd1,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd2,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd2}};

parameter bit [1:0] SpriteTableB_2_23[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd2,2'd3,2'd3},
'{2'd2,2'd3,2'd2,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2},
'{2'd3,2'd2,2'd2,2'd2,2'd2,2'd1,2'd3,2'd3},
'{2'd2,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_2_24[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_2_25[7:0][7:0] = '{'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_2_26[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_2_27[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_2_28[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd1,2'd1,2'd1,2'd3,2'd1,2'd3,2'd3,2'd2},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_2_29[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd2,2'd1,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd2,2'd1},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_2_30[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_2_31[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_2_32[7:0][7:0] = '{'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd1,2'd1,2'd3},
'{2'd2,2'd3,2'd1,2'd1,2'd1,2'd1,2'd1,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_2_33[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2}};

parameter bit [1:0] SpriteTableB_2_34[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_2_35[7:0][7:0] = '{'{2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_3_0[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_3_1[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_3_2[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_3_3[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2}};

parameter bit [1:0] SpriteTableB_3_4[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_3_5[7:0][7:0] = '{'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_3_6[7:0][7:0] = '{'{2'd1,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd1},
'{2'd1,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3,2'd1},
'{2'd1,2'd1,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_3_7[7:0][7:0] = '{'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd1,2'd1},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_3_8[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2},
'{2'd1,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2},
'{2'd1,2'd3,2'd2,2'd3,2'd3,2'd1,2'd2,2'd2},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd1,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_3_9[7:0][7:0] = '{'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd2,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_3_10[7:0][7:0] = '{'{2'd1,2'd1,2'd2,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd1,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_3_11[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_3_12[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd2,2'd2,2'd1,2'd1,2'd2,2'd1,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_3_13[7:0][7:0] = '{'{2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd3,2'd3},
'{2'd3,2'd1,2'd2,2'd2,2'd2,2'd1,2'd3,2'd3},
'{2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1},
'{2'd1,2'd1,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd2,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_3_14[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_3_15[7:0][7:0] = '{'{2'd3,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd2,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3}};

parameter bit [1:0] SpriteTableB_3_16[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_3_17[7:0][7:0] = '{'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3}};

parameter bit [1:0] SpriteTableB_3_18[7:0][7:0] = '{'{2'd2,2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_3_19[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd2,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_3_20[7:0][7:0] = '{'{2'd3,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_3_21[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_3_22[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_3_23[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd2,2'd2,2'd2,2'd1},
'{2'd2,2'd1,2'd1,2'd3,2'd1,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_3_24[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd1,2'd3,2'd1,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd2},
'{2'd1,2'd1,2'd3,2'd3,2'd2,2'd3,2'd2,2'd2},
'{2'd3,2'd1,2'd3,2'd1,2'd1,2'd3,2'd2,2'd2}};

parameter bit [1:0] SpriteTableB_3_25[7:0][7:0] = '{'{2'd3,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1},
'{2'd3,2'd3,2'd1,2'd2,2'd2,2'd1,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd3,2'd2,2'd2,2'd2,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd2,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd1,2'd3,2'd3,2'd2,2'd2,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_3_26[7:0][7:0] = '{'{2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_3_27[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_3_28[7:0][7:0] = '{'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_3_29[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_3_30[7:0][7:0] = '{'{2'd3,2'd3,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1}};

parameter bit [1:0] SpriteTableB_3_31[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_3_32[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd1,2'd2},
'{2'd3,2'd1,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_3_33[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd2,2'd2,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_3_34[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_3_35[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_4_0[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_4_1[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_4_2[7:0][7:0] = '{'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_4_3[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_4_4[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1}};

parameter bit [1:0] SpriteTableB_4_5[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_4_6[7:0][7:0] = '{'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd1,2'd3,2'd3,2'd1,2'd1,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_4_7[7:0][7:0] = '{'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_4_8[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd2,2'd1,2'd3,2'd3,2'd3},
'{2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_4_9[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd2,2'd2,2'd3,2'd3},
'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd2,2'd1,2'd1,2'd2,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_4_10[7:0][7:0] = '{'{2'd3,2'd1,2'd2,2'd2,2'd2,2'd1,2'd3,2'd3},
'{2'd1,2'd2,2'd2,2'd1,2'd1,2'd1,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd3,2'd2},
'{2'd3,2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd3},
'{2'd3,2'd3,2'd1,2'd1,2'd2,2'd2,2'd2,2'd3},
'{2'd3,2'd3,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd1,2'd2,2'd3,2'd3,2'd2}};

parameter bit [1:0] SpriteTableB_4_11[7:0][7:0] = '{'{2'd3,2'd3,2'd1,2'd2,2'd2,2'd2,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2}};

parameter bit [1:0] SpriteTableB_4_12[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_4_13[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd1,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd2},
'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd2,2'd2,2'd3}};

parameter bit [1:0] SpriteTableB_4_14[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_4_15[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_4_16[7:0][7:0] = '{'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_4_17[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_4_18[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_4_19[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_4_20[7:0][7:0] = '{'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_4_21[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_4_22[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_4_23[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd1,2'd3,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_4_24[7:0][7:0] = '{'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd1},
'{2'd3,2'd2,2'd1,2'd3,2'd3,2'd1,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_4_25[7:0][7:0] = '{'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd2},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd1,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2}};

parameter bit [1:0] SpriteTableB_4_26[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd3,2'd1,2'd1},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd1,2'd3,2'd3,2'd1,2'd1}};

parameter bit [1:0] SpriteTableB_4_27[7:0][7:0] = '{'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd2,2'd3,2'd1,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_4_28[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd1,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2}};

parameter bit [1:0] SpriteTableB_4_29[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_4_30[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_4_31[7:0][7:0] = '{'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_4_32[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd2,2'd1,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_4_33[7:0][7:0] = '{'{2'd3,2'd2,2'd1,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_4_34[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_4_35[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_5_0[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_5_1[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_5_2[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd1,2'd2,2'd2,2'd2,2'd2}};

parameter bit [1:0] SpriteTableB_5_3[7:0][7:0] = '{'{2'd3,2'd3,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_5_4[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd2,2'd3}};

parameter bit [1:0] SpriteTableB_5_5[7:0][7:0] = '{'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd1,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_5_6[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd2,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd1,2'd2,2'd2,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_5_7[7:0][7:0] = '{'{2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_5_8[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd2,2'd1,2'd2,2'd1,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_5_9[7:0][7:0] = '{'{2'd3,2'd3,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_5_10[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd1,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_5_11[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd2,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3},
'{2'd2,2'd2,2'd2,2'd3,2'd2,2'd2,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_5_12[7:0][7:0] = '{'{2'd2,2'd2,2'd3,2'd2,2'd2,2'd2,2'd1,2'd3},
'{2'd2,2'd2,2'd3,2'd2,2'd2,2'd2,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd2,2'd3,2'd2,2'd2,2'd3,2'd2,2'd3,2'd3},
'{2'd2,2'd3,2'd2,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd2,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd1,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_5_13[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_5_14[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_5_15[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_5_16[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_5_17[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_5_18[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_5_19[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_5_20[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_5_21[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_5_22[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd3}};

parameter bit [1:0] SpriteTableB_5_23[7:0][7:0] = '{'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd2,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd1,2'd3},
'{2'd3,2'd3,2'd2,2'd2,2'd2,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd2,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_5_24[7:0][7:0] = '{'{2'd1,2'd1,2'd2,2'd3,2'd2,2'd3,2'd1,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd2,2'd3,2'd2,2'd3},
'{2'd1,2'd2,2'd3,2'd3,2'd2,2'd3,2'd2,2'd3},
'{2'd3,2'd2,2'd2,2'd3,2'd2,2'd3,2'd2,2'd3},
'{2'd3,2'd1,2'd2,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd1,2'd2,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd1},
'{2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd2}};

parameter bit [1:0] SpriteTableB_5_25[7:0][7:0] = '{'{2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2},
'{2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd1,2'd2,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2},
'{2'd1,2'd2,2'd3,2'd3,2'd2,2'd2,2'd2,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3},
'{2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3},
'{2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3},
'{2'd2,2'd3,2'd2,2'd2,2'd2,2'd3,2'd3,2'd2}};

parameter bit [1:0] SpriteTableB_5_26[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd3},
'{2'd3,2'd3,2'd2,2'd2,2'd1,2'd3,2'd1,2'd3},
'{2'd2,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd1},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd2,2'd1,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd1,2'd2,2'd2,2'd2,2'd1,2'd3,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_5_27[7:0][7:0] = '{'{2'd2,2'd2,2'd1,2'd2,2'd2,2'd1,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd1,2'd1,2'd3,2'd3,2'd1},
'{2'd2,2'd2,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd1,2'd3},
'{2'd2,2'd1,2'd1,2'd1,2'd2,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_5_28[7:0][7:0] = '{'{2'd1,2'd2,2'd2,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd2,2'd1,2'd3,2'd1,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd2,2'd1,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_5_29[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd2,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_5_30[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_5_31[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_5_32[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_5_33[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_5_34[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_5_35[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_6_0[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd2,2'd1,2'd1,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_6_1[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_6_2[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_6_3[7:0][7:0] = '{'{2'd1,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd2,2'd3,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd2,2'd2,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2}};

parameter bit [1:0] SpriteTableB_6_4[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_6_5[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd1},
'{2'd2,2'd3,2'd3,2'd2,2'd2,2'd2,2'd3,2'd1},
'{2'd3,2'd1,2'd3,2'd2,2'd2,2'd2,2'd1,2'd2},
'{2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1},
'{2'd3,2'd1,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_6_6[7:0][7:0] = '{'{2'd3,2'd1,2'd3,2'd3,2'd1,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_6_7[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd1,2'd3,2'd1,2'd3,2'd1},
'{2'd2,2'd2,2'd2,2'd1,2'd3,2'd1,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd1,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd1,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_6_8[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_6_9[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd1,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_6_10[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd2,2'd2,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd2},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd2}};

parameter bit [1:0] SpriteTableB_6_11[7:0][7:0] = '{'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd1,2'd3,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd1,2'd3,2'd2,2'd2,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd2,2'd2,2'd3,2'd2,2'd2},
'{2'd3,2'd1,2'd3,2'd3,2'd2,2'd3,2'd3,2'd2}};

parameter bit [1:0] SpriteTableB_6_12[7:0][7:0] = '{'{2'd3,2'd1,2'd3,2'd2,2'd2,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_6_13[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_6_14[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_6_15[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd1,2'd3,2'd3,2'd2,2'd3}};

parameter bit [1:0] SpriteTableB_6_16[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_6_17[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_6_18[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_6_19[7:0][7:0] = '{'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_6_20[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_6_21[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd1,2'd3,2'd3,2'd1,2'd3,2'd3,2'd2,2'd3},
'{2'd1,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_6_22[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_6_23[7:0][7:0] = '{'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_6_24[7:0][7:0] = '{'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd2,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_6_25[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd2,2'd1,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd2,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_6_26[7:0][7:0] = '{'{2'd1,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd1},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_6_27[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd2,2'd2,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_6_28[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_6_29[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd2},
'{2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2}};

parameter bit [1:0] SpriteTableB_6_30[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_6_31[7:0][7:0] = '{'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_6_32[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_6_33[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_6_34[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_6_35[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_7_0[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_7_1[7:0][7:0] = '{'{2'd2,2'd2,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_7_2[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_7_3[7:0][7:0] = '{'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd1,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_7_4[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_7_5[7:0][7:0] = '{'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd1,2'd3,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_7_6[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_7_7[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_7_8[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd2}};

parameter bit [1:0] SpriteTableB_7_9[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd1,2'd3,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd3,2'd2},
'{2'd1,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd2,2'd3,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd2,2'd2,2'd3,2'd2,2'd2,2'd3,2'd2},
'{2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2}};

parameter bit [1:0] SpriteTableB_7_10[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd3,2'd3,2'd2,2'd3,2'd3,2'd2},
'{2'd2,2'd2,2'd3,2'd3,2'd2,2'd2,2'd3,2'd2},
'{2'd2,2'd2,2'd3,2'd2,2'd2,2'd2,2'd2,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd3,2'd2,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_7_11[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd2,2'd2,2'd2,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd2,2'd2,2'd2,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd2,2'd3,2'd2,2'd2,2'd3,2'd2,2'd3},
'{2'd3,2'd2,2'd2,2'd3,2'd2,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_7_12[7:0][7:0] = '{'{2'd3,2'd2,2'd2,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_7_13[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_7_14[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_7_15[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_7_16[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_7_17[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_7_18[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_7_19[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_7_20[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_7_21[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_7_22[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_7_23[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_7_24[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_7_25[7:0][7:0] = '{'{2'd2,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_7_26[7:0][7:0] = '{'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd1,2'd3,2'd1,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd1,2'd3,2'd1,2'd1}};

parameter bit [1:0] SpriteTableB_7_27[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd1,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd2,2'd2,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd1}};

parameter bit [1:0] SpriteTableB_7_28[7:0][7:0] = '{'{2'd3,2'd1,2'd3,2'd1,2'd3,2'd3,2'd2,2'd1},
'{2'd1,2'd3,2'd3,2'd3,2'd2,2'd3,2'd2,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd1,2'd2},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd3,2'd1},
'{2'd3,2'd3,2'd1,2'd2,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd1,2'd2,2'd2,2'd1,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_7_29[7:0][7:0] = '{'{2'd1,2'd2,2'd2,2'd2,2'd1,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd1,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd3,2'd1},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd1},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_7_30[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd1},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd1,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd3,2'd1,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_7_31[7:0][7:0] = '{'{2'd1,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd2,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_7_32[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_7_33[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_7_34[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_7_35[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_8_0[7:0][7:0] = '{'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_8_1[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_8_2[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd2,2'd2}};

parameter bit [1:0] SpriteTableB_8_3[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd2,2'd1,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_8_4[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_8_5[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd1,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_8_6[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_8_7[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_8_8[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2},
'{2'd1,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd2,2'd2,2'd2,2'd3,2'd2,2'd2,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd3,2'd2,2'd2,2'd3,2'd2,2'd2,2'd3}};

parameter bit [1:0] SpriteTableB_8_9[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd3,2'd2,2'd2,2'd3,2'd2,2'd2,2'd3},
'{2'd2,2'd3,2'd2,2'd2,2'd3,2'd2,2'd2,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3},
'{2'd2,2'd3,2'd2,2'd2,2'd3,2'd2,2'd3,2'd1},
'{2'd2,2'd3,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_8_10[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd1,2'd3},
'{2'd2,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd2,2'd2,2'd3,2'd1,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd2,2'd3,2'd1,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_8_11[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_8_12[7:0][7:0] = '{'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_8_13[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_8_14[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_8_15[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_8_16[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_8_17[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2}};

parameter bit [1:0] SpriteTableB_8_18[7:0][7:0] = '{'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd2,2'd3,2'd3,2'd2,2'd2,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd2,2'd2,2'd2},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_8_19[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_8_20[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_8_21[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_8_22[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_8_23[7:0][7:0] = '{'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_8_24[7:0][7:0] = '{'{2'd3,2'd3,2'd1,2'd1,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_8_25[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_8_26[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_8_27[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd1,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd1,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd1,2'd1,2'd2}};

parameter bit [1:0] SpriteTableB_8_28[7:0][7:0] = '{'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd1,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2},
'{2'd1,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_8_29[7:0][7:0] = '{'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_8_30[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_8_31[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_8_32[7:0][7:0] = '{'{2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_8_33[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_8_34[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_8_35[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_9_0[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3},
'{2'd3,2'd3,2'd1,2'd1,2'd1,2'd2,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_9_1[7:0][7:0] = '{'{2'd3,2'd3,2'd1,2'd2,2'd2,2'd2,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd1},
'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd1,2'd2,2'd2,2'd2,2'd2,2'd3},
'{2'd3,2'd3,2'd2,2'd1,2'd1,2'd2,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_9_2[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd2,2'd1,2'd3,2'd3,2'd3},
'{2'd2,2'd1,2'd1,2'd2,2'd2,2'd1,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_9_3[7:0][7:0] = '{'{2'd3,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd3},
'{2'd3,2'd3,2'd2,2'd2,2'd2,2'd1,2'd3,2'd3},
'{2'd1,2'd3,2'd2,2'd1,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd1,2'd2,2'd1,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_9_4[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_9_5[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_9_6[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1}};

parameter bit [1:0] SpriteTableB_9_7[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2}};

parameter bit [1:0] SpriteTableB_9_8[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd3,2'd2,2'd2,2'd3,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd3,2'd2,2'd2,2'd3,2'd2,2'd2}};

parameter bit [1:0] SpriteTableB_9_9[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd2,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_9_10[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd2,2'd3}};

parameter bit [1:0] SpriteTableB_9_11[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_9_12[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_9_13[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_9_14[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_9_15[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_9_16[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_9_17[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd2,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd1,2'd1,2'd2},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3}};

parameter bit [1:0] SpriteTableB_9_18[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd3,2'd3,2'd2,2'd2,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd2,2'd2,2'd3},
'{2'd3,2'd2,2'd2,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd2,2'd1,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_9_19[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_9_20[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_9_21[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_9_22[7:0][7:0] = '{'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_9_23[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_9_24[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_9_25[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_9_26[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd2,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_9_27[7:0][7:0] = '{'{2'd3,2'd2,2'd2,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd2,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd2,2'd2,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd2,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd2},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_9_28[7:0][7:0] = '{'{2'd3,2'd3,2'd2,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_9_29[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_9_30[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_9_31[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_9_32[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd2,2'd1},
'{2'd2,2'd1,2'd1,2'd1,2'd2,2'd3,2'd2,2'd1}};

parameter bit [1:0] SpriteTableB_9_33[7:0][7:0] = '{'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd1,2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd2},
'{2'd1,2'd2,2'd3,2'd3,2'd3,2'd2,2'd3,2'd2}};

parameter bit [1:0] SpriteTableB_9_34[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_9_35[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_10_0[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_10_1[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_10_2[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_10_3[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_10_4[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd1,2'd1,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd1,2'd2,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd2,2'd3},
'{2'd3,2'd1,2'd3,2'd1,2'd2,2'd2,2'd2,2'd2}};

parameter bit [1:0] SpriteTableB_10_5[7:0][7:0] = '{'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_10_6[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_10_7[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3}};

parameter bit [1:0] SpriteTableB_10_8[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd2,2'd2,2'd3,2'd2,2'd2,2'd3,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd2,2'd2,2'd3,2'd2,2'd2,2'd3,2'd2}};

parameter bit [1:0] SpriteTableB_10_9[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd2,2'd2,2'd3,2'd2,2'd2,2'd3,2'd2},
'{2'd3,2'd3,2'd2,2'd3,2'd2,2'd2,2'd3,2'd2},
'{2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd1,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1}};

parameter bit [1:0] SpriteTableB_10_10[7:0][7:0] = '{'{2'd3,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_10_11[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_10_12[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_10_13[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_10_14[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_10_15[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_10_16[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_10_17[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd2}};

parameter bit [1:0] SpriteTableB_10_18[7:0][7:0] = '{'{2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd2},
'{2'd2,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_10_19[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_10_20[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_10_21[7:0][7:0] = '{'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_10_22[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_10_23[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_10_24[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_10_25[7:0][7:0] = '{'{2'd1,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_10_26[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_10_27[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1},
'{2'd2,2'd1,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd1},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd1,2'd1}};

parameter bit [1:0] SpriteTableB_10_28[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd1,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd1,2'd1,2'd3},
'{2'd3,2'd3,2'd1,2'd1,2'd1,2'd1,2'd1,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd1,2'd1,2'd1,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd1,2'd3},
'{2'd3,2'd1,2'd1,2'd3,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd1,2'd1,2'd1,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_10_29[7:0][7:0] = '{'{2'd3,2'd1,2'd3,2'd1,2'd1,2'd1,2'd3,2'd1},
'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_10_30[7:0][7:0] = '{'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_10_31[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_10_32[7:0][7:0] = '{'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1},
'{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_10_33[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_10_34[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_10_35[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_11_0[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd2,2'd1,2'd1,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_11_1[7:0][7:0] = '{'{2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd2},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2}};

parameter bit [1:0] SpriteTableB_11_2[7:0][7:0] = '{'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1},
'{2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_11_3[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_11_4[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd2,2'd2,2'd2,2'd2,2'd3}};

parameter bit [1:0] SpriteTableB_11_5[7:0][7:0] = '{'{2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_11_6[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1}};

parameter bit [1:0] SpriteTableB_11_7[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_11_8[7:0][7:0] = '{'{2'd2,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd3,2'd1,2'd3,2'd3,2'd1},
'{2'd2,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd3,2'd1,2'd3,2'd3},
'{2'd2,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_11_9[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd2,2'd2,2'd3,2'd3,2'd1,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_11_10[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd1},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_11_11[7:0][7:0] = '{'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_11_12[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_11_13[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_11_14[7:0][7:0] = '{'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_11_15[7:0][7:0] = '{'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_11_16[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_11_17[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd2,2'd3,2'd1,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_11_18[7:0][7:0] = '{'{2'd2,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd2,2'd2,2'd3,2'd3,2'd1,2'd3},
'{2'd2,2'd3,2'd3,2'd2,2'd3,2'd3,2'd1,2'd3},
'{2'd2,2'd3,2'd3,2'd2,2'd2,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_11_19[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_11_20[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_11_21[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_11_22[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_11_23[7:0][7:0] = '{'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_11_24[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd1,2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_11_25[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd1,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_11_26[7:0][7:0] = '{'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd1,2'd1,2'd3,2'd3,2'd1,2'd3,2'd2,2'd3},
'{2'd1,2'd1,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_11_27[7:0][7:0] = '{'{2'd1,2'd3,2'd3,2'd3,2'd2,2'd2,2'd3,2'd3},
'{2'd1,2'd3,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2},
'{2'd1,2'd3,2'd2,2'd1,2'd3,2'd3,2'd2,2'd2},
'{2'd1,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd1,2'd3,2'd3,2'd1,2'd1,2'd3,2'd1},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_11_28[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1},
'{2'd1,2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_11_29[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_11_30[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_11_31[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd1,2'd3,2'd1,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_11_32[7:0][7:0] = '{'{2'd3,2'd3,2'd1,2'd3,2'd1,2'd1,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd3},
'{2'd3,2'd1,2'd2,2'd1,2'd2,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd1,2'd2,2'd2,2'd3,2'd2,2'd2}};

parameter bit [1:0] SpriteTableB_11_33[7:0][7:0] = '{'{2'd3,2'd3,2'd2,2'd3,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd1,2'd2,2'd1,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_11_34[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_11_35[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_12_0[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_12_1[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd2,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd2,2'd2,2'd1,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_12_2[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd1,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_12_3[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_12_4[7:0][7:0] = '{'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd3},
'{2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_12_5[7:0][7:0] = '{'{2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd3},
'{2'd2,2'd3,2'd2,2'd2,2'd2,2'd3,2'd2,2'd3},
'{2'd2,2'd3,2'd2,2'd2,2'd2,2'd3,2'd3,2'd1},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2}};

parameter bit [1:0] SpriteTableB_12_6[7:0][7:0] = '{'{2'd2,2'd3,2'd2,2'd2,2'd2,2'd3,2'd2,2'd2},
'{2'd2,2'd3,2'd2,2'd2,2'd2,2'd3,2'd3,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1},
'{2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd3},
'{2'd2,2'd3,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd2,2'd2,2'd2,2'd3,2'd2,2'd3}};

parameter bit [1:0] SpriteTableB_12_7[7:0][7:0] = '{'{2'd3,2'd3,2'd1,2'd2,2'd2,2'd2,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd2,2'd2,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd1},
'{2'd1,2'd3,2'd1,2'd3,2'd3,2'd1,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_12_8[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd1,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd2},
'{2'd1,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd2}};

parameter bit [1:0] SpriteTableB_12_9[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd2,2'd2},
'{2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2}};

parameter bit [1:0] SpriteTableB_12_10[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd1,2'd3,2'd2,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd1,2'd3,2'd2,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd2},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_12_11[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_12_12[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_12_13[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_12_14[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_12_15[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_12_16[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_12_17[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd2,2'd2,2'd3,2'd2,2'd2},
'{2'd3,2'd1,2'd3,2'd2,2'd1,2'd1,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_12_18[7:0][7:0] = '{'{2'd3,2'd1,2'd3,2'd2,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd2,2'd1,2'd2,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd2,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd2,2'd2,2'd3,2'd2,2'd3},
'{2'd3,2'd1,2'd3,2'd2,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_12_19[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd3}};

parameter bit [1:0] SpriteTableB_12_20[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_12_21[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_12_22[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2},
'{2'd1,2'd2,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_12_23[7:0][7:0] = '{'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd2,2'd1,2'd2},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_12_24[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_12_25[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_12_26[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_12_27[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd3},
'{2'd2,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd2},
'{2'd2,2'd3,2'd2,2'd2,2'd2,2'd3,2'd2,2'd3},
'{2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd2}};

parameter bit [1:0] SpriteTableB_12_28[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd1},
'{2'd1,2'd3,2'd2,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd1,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_12_29[7:0][7:0] = '{'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd1},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd1,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_12_30[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd1},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_12_31[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd1,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_12_32[7:0][7:0] = '{'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd2},
'{2'd2,2'd3,2'd2,2'd3,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd2,2'd2,2'd3,2'd2,2'd2,2'd3},
'{2'd1,2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd2,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd2,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2}};

parameter bit [1:0] SpriteTableB_12_33[7:0][7:0] = '{'{2'd1,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_12_34[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_12_35[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_13_0[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_13_1[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_13_2[7:0][7:0] = '{'{2'd1,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_13_3[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_13_4[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_13_5[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd1,2'd1},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd1,2'd2},
'{2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd2,2'd2,2'd2,2'd1,2'd3,2'd3,2'd3,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_13_6[7:0][7:0] = '{'{2'd2,2'd2,2'd3,2'd2,2'd1,2'd3,2'd2,2'd3},
'{2'd2,2'd2,2'd3,2'd1,2'd3,2'd3,2'd2,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd1,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd1,2'd2,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_13_7[7:0][7:0] = '{'{2'd3,2'd1,2'd1,2'd2,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd2,2'd3,2'd2,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_13_8[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd2,2'd2,2'd3,2'd2,2'd2,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_13_9[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd2,2'd2,2'd3,2'd2,2'd2,2'd3,2'd2},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd2,2'd3,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd2,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3}};

parameter bit [1:0] SpriteTableB_13_10[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd2,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd2,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd1},
'{2'd3,2'd3,2'd2,2'd3,2'd2,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_13_11[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_13_12[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_13_13[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd2,2'd1,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_13_14[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_13_15[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_13_16[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd1,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd1,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_13_17[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_13_18[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_13_19[7:0][7:0] = '{'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_13_20[7:0][7:0] = '{'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_13_21[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd2,2'd3,2'd2,2'd3,2'd3,2'd3,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_13_22[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_13_23[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_13_24[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_13_25[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_13_26[7:0][7:0] = '{'{2'd3,2'd3,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_13_27[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd2,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_13_28[7:0][7:0] = '{'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd2,2'd3,2'd2,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd2},
'{2'd3,2'd1,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_13_29[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd2,2'd3,2'd2,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd2,2'd2,2'd2,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd2,2'd1,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2}};

parameter bit [1:0] SpriteTableB_13_30[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd1,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd1,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd1,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd2,2'd2}};

parameter bit [1:0] SpriteTableB_13_31[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd1,2'd2,2'd2,2'd2,2'd1},
'{2'd3,2'd1,2'd3,2'd1,2'd1,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd1,2'd3,2'd1,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_13_32[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd2,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_13_33[7:0][7:0] = '{'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd1},
'{2'd1,2'd2,2'd3,2'd3,2'd3,2'd1,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd1,2'd2},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd2}};

parameter bit [1:0] SpriteTableB_13_34[7:0][7:0] = '{'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_13_35[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_14_0[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1},
'{2'd3,2'd1,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_14_1[7:0][7:0] = '{'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_14_2[7:0][7:0] = '{'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_14_3[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd1,2'd3,2'd3,2'd1,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_14_4[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_14_5[7:0][7:0] = '{'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd1},
'{2'd2,2'd3,2'd2,2'd1,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd1,2'd2},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_14_6[7:0][7:0] = '{'{2'd3,2'd2,2'd3,2'd2,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd2,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_14_7[7:0][7:0] = '{'{2'd2,2'd3,2'd2,2'd2,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd1},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_14_8[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd3,2'd3,2'd2,2'd3,2'd3,2'd2,2'd3}};

parameter bit [1:0] SpriteTableB_14_9[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd1,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd1,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd1,2'd3,2'd2,2'd3,2'd3,2'd2,2'd3},
'{2'd1,2'd1,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2}};

parameter bit [1:0] SpriteTableB_14_10[7:0][7:0] = '{'{2'd1,2'd1,2'd3,2'd2,2'd2,2'd2,2'd3,2'd2},
'{2'd3,2'd1,2'd3,2'd2,2'd2,2'd3,2'd2,2'd3},
'{2'd3,2'd1,2'd3,2'd2,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd1,2'd3,2'd2,2'd3,2'd2,2'd2,2'd2},
'{2'd3,2'd1,2'd2,2'd2,2'd2,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd3}};

parameter bit [1:0] SpriteTableB_14_11[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd3},
'{2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3},
'{2'd1,2'd3,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd2,2'd3,2'd2,2'd3},
'{2'd1,2'd3,2'd3,2'd2,2'd3,2'd3,2'd2,2'd3}};

parameter bit [1:0] SpriteTableB_14_12[7:0][7:0] = '{'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_14_13[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_14_14[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_14_15[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_14_16[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_14_17[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_14_18[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_14_19[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_14_20[7:0][7:0] = '{'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_14_21[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_14_22[7:0][7:0] = '{'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_14_23[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd2,2'd1},
'{2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3}};

parameter bit [1:0] SpriteTableB_14_24[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_14_25[7:0][7:0] = '{'{2'd3,2'd2,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd2,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_14_26[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_14_27[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_14_28[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2}};

parameter bit [1:0] SpriteTableB_14_29[7:0][7:0] = '{'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd2,2'd3,2'd2},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd2,2'd3,2'd2}};

parameter bit [1:0] SpriteTableB_14_30[7:0][7:0] = '{'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd2,2'd2,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd2,2'd3},
'{2'd2,2'd3,2'd2,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd2,2'd3,2'd3,2'd2,2'd2,2'd3,2'd2,2'd3},
'{2'd1,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd2,2'd3,2'd2,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_14_31[7:0][7:0] = '{'{2'd3,2'd1,2'd3,2'd2,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd1},
'{2'd1,2'd3,2'd2,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd2,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_14_32[7:0][7:0] = '{'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_14_33[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_14_34[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_14_35[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_15_0[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_15_1[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_15_2[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_15_3[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd1},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd2,2'd2,2'd1},
'{2'd1,2'd1,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2}};

parameter bit [1:0] SpriteTableB_15_4[7:0][7:0] = '{'{2'd3,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd1,2'd3,2'd1},
'{2'd3,2'd3,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_15_5[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_15_6[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd2,2'd1,2'd2,2'd1,2'd3,2'd3},
'{2'd3,2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1},
'{2'd3,2'd3,2'd2,2'd2,2'd1,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd3}};

parameter bit [1:0] SpriteTableB_15_7[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd1,2'd1,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1},
'{2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_15_8[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd1},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd1},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd1},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd1},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd1},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd1},
'{2'd3,2'd2,2'd3,2'd3,2'd2,2'd2,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_15_9[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd1},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3},
'{2'd3,2'd2,2'd2,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd2,2'd3,2'd2,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_15_10[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd1,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd1,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd2,2'd3,2'd1,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd2,2'd3,2'd1,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd2,2'd3,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_15_11[7:0][7:0] = '{'{2'd2,2'd2,2'd3,2'd3,2'd2,2'd3,2'd1,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd1,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd1,2'd3},
'{2'd3,2'd2,2'd2,2'd1,2'd2,2'd3,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_15_12[7:0][7:0] = '{'{2'd3,2'd2,2'd3,2'd2,2'd2,2'd3,2'd1,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_15_13[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_15_14[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_15_15[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_15_16[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_15_17[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_15_18[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_15_19[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_15_20[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_15_21[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_15_22[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_15_23[7:0][7:0] = '{'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd1,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_15_24[7:0][7:0] = '{'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_15_25[7:0][7:0] = '{'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd1,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd1,2'd2,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_15_26[7:0][7:0] = '{'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_15_27[7:0][7:0] = '{'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd2,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd2,2'd1,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_15_28[7:0][7:0] = '{'{2'd3,2'd1,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd2,2'd3,2'd2,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2}};

parameter bit [1:0] SpriteTableB_15_29[7:0][7:0] = '{'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd2,2'd2},
'{2'd2,2'd1,2'd2,2'd3,2'd3,2'd3,2'd2,2'd2},
'{2'd2,2'd3,2'd1,2'd3,2'd3,2'd1,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_15_30[7:0][7:0] = '{'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_15_31[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_15_32[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_15_33[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_15_34[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_15_35[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_16_0[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_16_1[7:0][7:0] = '{'{2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_16_2[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_16_3[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd1,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_16_4[7:0][7:0] = '{'{2'd2,2'd1,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd2,2'd1,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd2,2'd1,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd2,2'd1,2'd1,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd1,2'd1,2'd3,2'd1},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd1,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_16_5[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1}};

parameter bit [1:0] SpriteTableB_16_6[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd1,2'd2,2'd2,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd1,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd1,2'd3,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_16_7[7:0][7:0] = '{'{2'd2,2'd2,2'd1,2'd2,2'd3,2'd2,2'd1,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_16_8[7:0][7:0] = '{'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_16_9[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_16_10[7:0][7:0] = '{'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3,2'd1},
'{2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd1,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_16_11[7:0][7:0] = '{'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd1,2'd3,2'd2},
'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd2}};

parameter bit [1:0] SpriteTableB_16_12[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_16_13[7:0][7:0] = '{'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_16_14[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_16_15[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_16_16[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_16_17[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_16_18[7:0][7:0] = '{'{2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_16_19[7:0][7:0] = '{'{2'd1,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_16_20[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_16_21[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_16_22[7:0][7:0] = '{'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_16_23[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_16_24[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_16_25[7:0][7:0] = '{'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd2,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd2,2'd2,2'd3},
'{2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd2,2'd2},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_16_26[7:0][7:0] = '{'{2'd3,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_16_27[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2}};

parameter bit [1:0] SpriteTableB_16_28[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_16_29[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd3,2'd2,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd1,2'd1,2'd2,2'd3,2'd2,2'd2,2'd2},
'{2'd1,2'd1,2'd3,2'd3,2'd2,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd2}};

parameter bit [1:0] SpriteTableB_16_30[7:0][7:0] = '{'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_16_31[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_16_32[7:0][7:0] = '{'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3}};

parameter bit [1:0] SpriteTableB_16_33[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_16_34[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_16_35[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_17_0[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_17_1[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_17_2[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd2,2'd2,2'd2,2'd1,2'd3,2'd3,2'd1,2'd2},
'{2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2}};

parameter bit [1:0] SpriteTableB_17_3[7:0][7:0] = '{'{2'd3,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd3,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd2,2'd2,2'd3,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd2,2'd2,2'd3,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd2,2'd2,2'd3,2'd3,2'd1,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2}};

parameter bit [1:0] SpriteTableB_17_4[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd2,2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd1},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_17_5[7:0][7:0] = '{'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd1,2'd1,2'd1,2'd3,2'd1},
'{2'd1,2'd3,2'd3,2'd1,2'd3,2'd1,2'd3,2'd1},
'{2'd1,2'd3,2'd1,2'd1,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_17_6[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd1,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd1,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_17_7[7:0][7:0] = '{'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd1,2'd3,2'd3,2'd3,2'd1,2'd1},
'{2'd2,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd1}};

parameter bit [1:0] SpriteTableB_17_8[7:0][7:0] = '{'{2'd1,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd1,2'd3,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd1,2'd3,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd2,2'd2}};

parameter bit [1:0] SpriteTableB_17_9[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd1,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd1,2'd3,2'd2,2'd2,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd1,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd1,2'd3,2'd3,2'd2,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3}};

parameter bit [1:0] SpriteTableB_17_10[7:0][7:0] = '{'{2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd2,2'd2,2'd2,2'd3},
'{2'd2,2'd2,2'd2,2'd3,2'd2,2'd2,2'd2,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2},
'{2'd2,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd1,2'd2}};

parameter bit [1:0] SpriteTableB_17_11[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd3,2'd2,2'd2,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd2,2'd2,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2}};

parameter bit [1:0] SpriteTableB_17_12[7:0][7:0] = '{'{2'd3,2'd2,2'd3,2'd3,2'd2,2'd3,2'd2,2'd3},
'{2'd2,2'd3,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_17_13[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_17_14[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd1},
'{2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_17_15[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_17_16[7:0][7:0] = '{'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_17_17[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_17_18[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_17_19[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_17_20[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_17_21[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_17_22[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_17_23[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_17_24[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_17_25[7:0][7:0] = '{'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1},
'{2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_17_26[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1},
'{2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_17_27[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_17_28[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_17_29[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd3,2'd3,2'd2,2'd2,2'd2,2'd3,2'd2},
'{2'd2,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd2},
'{2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd1,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_17_30[7:0][7:0] = '{'{2'd1,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd1,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_17_31[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd1,2'd3,2'd1},
'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_17_32[7:0][7:0] = '{'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd1,2'd1,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd1,2'd3,2'd1,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_17_33[7:0][7:0] = '{'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_17_34[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_17_35[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_18_0[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_18_1[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_18_2[7:0][7:0] = '{'{2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd1,2'd2,2'd1,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd2,2'd3,2'd3,2'd1,2'd3},
'{2'd2,2'd2,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd2}};

parameter bit [1:0] SpriteTableB_18_3[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd3,2'd2,2'd2,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd3,2'd2,2'd2,2'd2,2'd3},
'{2'd2,2'd2,2'd3,2'd2,2'd2,2'd3,2'd3,2'd2},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd2,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2}};

parameter bit [1:0] SpriteTableB_18_4[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd1,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_18_5[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_18_6[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd1,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_18_7[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd1,2'd1,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd2,2'd2,2'd2,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_18_8[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd2,2'd2,2'd3,2'd2,2'd2,2'd3,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd2,2'd2,2'd3,2'd2,2'd2,2'd3,2'd2}};

parameter bit [1:0] SpriteTableB_18_9[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd2,2'd2,2'd3,2'd2,2'd2,2'd3,2'd2},
'{2'd3,2'd2,2'd2,2'd3,2'd2,2'd2,2'd3,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd2,2'd3,2'd3,2'd2,2'd3,2'd3,2'd2},
'{2'd3,2'd2,2'd2,2'd3,2'd2,2'd2,2'd3,2'd2}};

parameter bit [1:0] SpriteTableB_18_10[7:0][7:0] = '{'{2'd2,2'd3,2'd2,2'd2,2'd3,2'd2,2'd2,2'd2},
'{2'd3,2'd2,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd2,2'd3,2'd3,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd2,2'd3},
'{2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_18_11[7:0][7:0] = '{'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_18_12[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_18_13[7:0][7:0] = '{'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_18_14[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd1,2'd2,2'd2,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd1,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_18_15[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_18_16[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_18_17[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2}};

parameter bit [1:0] SpriteTableB_18_18[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_18_19[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_18_20[7:0][7:0] = '{'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd1,2'd3,2'd1,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_18_21[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_18_22[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_18_23[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_18_24[7:0][7:0] = '{'{2'd1,2'd3,2'd3,2'd1,2'd1,2'd1,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_18_25[7:0][7:0] = '{'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd1,2'd1,2'd1,2'd3,2'd1,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_18_26[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd1,2'd2},
'{2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd2,2'd2,2'd3}};

parameter bit [1:0] SpriteTableB_18_27[7:0][7:0] = '{'{2'd3,2'd1,2'd3,2'd3,2'd2,2'd2,2'd2,2'd3},
'{2'd1,2'd2,2'd3,2'd3,2'd2,2'd2,2'd2,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd2,2'd2,2'd2,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_18_28[7:0][7:0] = '{'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd2,2'd2,2'd2,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd3,2'd3,2'd2,2'd2,2'd2,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd2,2'd2,2'd2,2'd3}};

parameter bit [1:0] SpriteTableB_18_29[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd3,2'd2,2'd1,2'd1,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd1,2'd3,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_18_30[7:0][7:0] = '{'{2'd2,2'd2,2'd3,2'd3,2'd1,2'd3,2'd1,2'd3},
'{2'd2,2'd2,2'd2,2'd1,2'd3,2'd3,2'd3,2'd1},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_18_31[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_18_32[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_18_33[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd1,2'd1,2'd2,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_18_34[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd1,2'd1,2'd2,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_18_35[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_19_0[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_19_1[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_19_2[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_19_3[7:0][7:0] = '{'{2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd2,2'd2,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1},
'{2'd2,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_19_4[7:0][7:0] = '{'{2'd2,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd1,2'd2,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd2,2'd2,2'd2,2'd1,2'd1,2'd3},
'{2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd1,2'd1,2'd2,2'd3,2'd3,2'd2,2'd1,2'd2},
'{2'd1,2'd1,2'd2,2'd3,2'd3,2'd2,2'd2,2'd2}};

parameter bit [1:0] SpriteTableB_19_5[7:0][7:0] = '{'{2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd1,2'd2,2'd3,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd2,2'd2,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd1,2'd3,2'd1,2'd2,2'd3,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2}};

parameter bit [1:0] SpriteTableB_19_6[7:0][7:0] = '{'{2'd3,2'd1,2'd2,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd2,2'd2,2'd3,2'd3,2'd2,2'd3,2'd2},
'{2'd3,2'd2,2'd2,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd2,2'd2,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2}};

parameter bit [1:0] SpriteTableB_19_7[7:0][7:0] = '{'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_19_8[7:0][7:0] = '{'{2'd2,2'd3,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd1,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd1,2'd3},
'{2'd2,2'd3,2'd2,2'd2,2'd3,2'd3,2'd1,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd1,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_19_9[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd2,2'd2,2'd3,2'd1,2'd3,2'd3},
'{2'd2,2'd3,2'd2,2'd2,2'd3,2'd1,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd3,2'd1,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_19_10[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd2,2'd3,2'd1,2'd3,2'd3,2'd1},
'{2'd2,2'd3,2'd2,2'd3,2'd1,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_19_11[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_19_12[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd3}};

parameter bit [1:0] SpriteTableB_19_13[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_19_14[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_19_15[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_19_16[7:0][7:0] = '{'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_19_17[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd3},
'{2'd2,2'd3,2'd3,2'd2,2'd2,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd1},
'{2'd2,2'd3,2'd3,2'd3,2'd2,2'd2,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_19_18[7:0][7:0] = '{'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd2,2'd2,2'd2,2'd3,2'd1,2'd3},
'{2'd2,2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_19_19[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_19_20[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_19_21[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_19_22[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_19_23[7:0][7:0] = '{'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_19_24[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_19_25[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1}};

parameter bit [1:0] SpriteTableB_19_26[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3}};

parameter bit [1:0] SpriteTableB_19_27[7:0][7:0] = '{'{2'd3,2'd2,2'd2,2'd2,2'd3,2'd3,2'd2,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd2,2'd3,2'd2,2'd3},
'{2'd3,2'd2,2'd2,2'd3,2'd3,2'd2,2'd2,2'd3},
'{2'd3,2'd1,2'd2,2'd2,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd1,2'd1,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd1,2'd3,2'd1,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd2}};

parameter bit [1:0] SpriteTableB_19_28[7:0][7:0] = '{'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd2,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd2,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd2,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd2,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_19_29[7:0][7:0] = '{'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd1,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd1},
'{2'd1,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd1,2'd1,2'd2}};

parameter bit [1:0] SpriteTableB_19_30[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd2},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_19_31[7:0][7:0] = '{'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_19_32[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_19_33[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_19_34[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_19_35[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_20_0[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_20_1[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd1,2'd2,2'd2,2'd2,2'd2}};

parameter bit [1:0] SpriteTableB_20_2[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd1,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_20_3[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd1}};

parameter bit [1:0] SpriteTableB_20_4[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd2},
'{2'd3,2'd1,2'd3,2'd3,2'd2,2'd2,2'd1,2'd2},
'{2'd1,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd1,2'd2,2'd2,2'd2,2'd1},
'{2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd2,2'd3}};

parameter bit [1:0] SpriteTableB_20_5[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd2,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd2,2'd3,2'd2,2'd3,2'd2},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd2,2'd3,2'd2,2'd3,2'd2,2'd2,2'd2},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_20_6[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_20_7[7:0][7:0] = '{'{2'd2,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_20_8[7:0][7:0] = '{'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd1,2'd3,2'd2},
'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd2,2'd2}};

parameter bit [1:0] SpriteTableB_20_9[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd1,2'd3,2'd2,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd2,2'd2},
'{2'd3,2'd1,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd1,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd3,2'd2,2'd2},
'{2'd1,2'd3,2'd3,2'd2,2'd2,2'd3,2'd2,2'd2}};

parameter bit [1:0] SpriteTableB_20_10[7:0][7:0] = '{'{2'd1,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd2},
'{2'd3,2'd2,2'd2,2'd3,2'd3,2'd2,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_20_11[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_20_12[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_20_13[7:0][7:0] = '{'{2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_20_14[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_20_15[7:0][7:0] = '{'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_20_16[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_20_17[7:0][7:0] = '{'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_20_18[7:0][7:0] = '{'{2'd1,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd2},
'{2'd1,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_20_19[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_20_20[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_20_21[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_20_22[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_20_23[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_20_24[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_20_25[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_20_26[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd1,2'd3,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_20_27[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd1,2'd1,2'd1},
'{2'd2,2'd2,2'd3,2'd3,2'd1,2'd1,2'd3,2'd1},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd1,2'd3,2'd1},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd2,2'd3,2'd2,2'd3,2'd3,2'd3,2'd2,2'd2}};

parameter bit [1:0] SpriteTableB_20_28[7:0][7:0] = '{'{2'd3,2'd2,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd1,2'd1,2'd3,2'd1,2'd2,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_20_29[7:0][7:0] = '{'{2'd3,2'd1,2'd3,2'd3,2'd1,2'd2,2'd1,2'd2},
'{2'd1,2'd1,2'd3,2'd3,2'd1,2'd1,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd3},
'{2'd2,2'd3,2'd2,2'd2,2'd2,2'd1,2'd1,2'd3},
'{2'd3,2'd3,2'd2,2'd2,2'd1,2'd3,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_20_30[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd2,2'd1,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd2,2'd2,2'd2,2'd1,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd2,2'd1,2'd1,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_20_31[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_20_32[7:0][7:0] = '{'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_20_33[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_20_34[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd2}};

parameter bit [1:0] SpriteTableB_20_35[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd2,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_21_0[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_21_1[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd2,2'd1,2'd2,2'd2,2'd1,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd1,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd1,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_21_2[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_21_3[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1}};

parameter bit [1:0] SpriteTableB_21_4[7:0][7:0] = '{'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd3},
'{2'd2,2'd2,2'd1,2'd3,2'd2,2'd2,2'd2,2'd3},
'{2'd2,2'd2,2'd3,2'd2,2'd3,2'd3,2'd2,2'd3},
'{2'd2,2'd1,2'd2,2'd3,2'd2,2'd3,2'd2,2'd3},
'{2'd2,2'd2,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd3,2'd2,2'd2,2'd2,2'd2,2'd3},
'{2'd2,2'd2,2'd3,2'd2,2'd2,2'd2,2'd2,2'd3},
'{2'd2,2'd2,2'd3,2'd2,2'd2,2'd2,2'd2,2'd3}};

parameter bit [1:0] SpriteTableB_21_5[7:0][7:0] = '{'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3}};

parameter bit [1:0] SpriteTableB_21_6[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd2},
'{2'd1,2'd3,2'd3,2'd2,2'd3,2'd2,2'd3,2'd2},
'{2'd1,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_21_7[7:0][7:0] = '{'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd1,2'd3,2'd3,2'd2,2'd2,2'd1,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1},
'{2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2}};

parameter bit [1:0] SpriteTableB_21_8[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd2,2'd2,2'd3,2'd2,2'd2,2'd3,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd2,2'd2,2'd3,2'd2,2'd2,2'd3,2'd2}};

parameter bit [1:0] SpriteTableB_21_9[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd2,2'd2,2'd3,2'd2,2'd2,2'd3,2'd2},
'{2'd3,2'd2,2'd2,2'd3,2'd2,2'd2,2'd3,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd2,2'd2,2'd3,2'd2,2'd2,2'd3,2'd2},
'{2'd3,2'd2,2'd2,2'd3,2'd2,2'd2,2'd3,2'd3},
'{2'd3,2'd2,2'd2,2'd3,2'd2,2'd2,2'd3,2'd2}};

parameter bit [1:0] SpriteTableB_21_10[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd2,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_21_11[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_21_12[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_21_13[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_21_14[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_21_15[7:0][7:0] = '{'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_21_16[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd1},
'{2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_21_17[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_21_18[7:0][7:0] = '{'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd2,2'd2,2'd3,2'd3},
'{2'd3,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_21_19[7:0][7:0] = '{'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_21_20[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_21_21[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_21_22[7:0][7:0] = '{'{2'd3,2'd3,2'd2,2'd1,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_21_23[7:0][7:0] = '{'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_21_24[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd2},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_21_25[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd1,2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3},
'{2'd1,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_21_26[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd1,2'd3,2'd3,2'd1,2'd1,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_21_27[7:0][7:0] = '{'{2'd2,2'd2,2'd3,2'd2,2'd2,2'd2,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3},
'{2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_21_28[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_21_29[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd2},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_21_30[7:0][7:0] = '{'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd1,2'd2},
'{2'd1,2'd3,2'd1,2'd3,2'd3,2'd3,2'd1,2'd2}};

parameter bit [1:0] SpriteTableB_21_31[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd1,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd1},
'{2'd1,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_21_32[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_21_33[7:0][7:0] = '{'{2'd2,2'd1,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd2,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2}};

parameter bit [1:0] SpriteTableB_21_34[7:0][7:0] = '{'{2'd1,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd2},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1}};

parameter bit [1:0] SpriteTableB_21_35[7:0][7:0] = '{'{2'd3,2'd2,2'd1,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_22_0[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_22_1[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_22_2[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_22_3[7:0][7:0] = '{'{2'd3,2'd2,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd2,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_22_4[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd1,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd2,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_22_5[7:0][7:0] = '{'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd1,2'd3,2'd3,2'd3,2'd1},
'{2'd2,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_22_6[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_22_7[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd1},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_22_8[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd1},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd1,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd1,2'd3},
'{2'd2,2'd3,2'd2,2'd2,2'd3,2'd3,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_22_9[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd1,2'd2,2'd3,2'd1,2'd3},
'{2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd1,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd3,2'd1,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd2,2'd3,2'd1,2'd3,2'd3},
'{2'd2,2'd3,2'd2,2'd2,2'd3,2'd1,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_22_10[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd2,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_22_11[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_22_12[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_22_13[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_22_14[7:0][7:0] = '{'{2'd3,2'd3,2'd1,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_22_15[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd1,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd1,2'd1,2'd1,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd1,2'd1,2'd1,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_22_16[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_22_17[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_22_18[7:0][7:0] = '{'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_22_19[7:0][7:0] = '{'{2'd1,2'd3,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_22_20[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_22_21[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_22_22[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_22_23[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_22_24[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_22_25[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_22_26[7:0][7:0] = '{'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_22_27[7:0][7:0] = '{'{2'd3,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_22_28[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_22_29[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd1,2'd1},
'{2'd3,2'd2,2'd2,2'd2,2'd3,2'd3,2'd1,2'd1},
'{2'd3,2'd1,2'd2,2'd3,2'd3,2'd2,2'd1,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd2,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_22_30[7:0][7:0] = '{'{2'd3,2'd3,2'd1,2'd3,2'd2,2'd2,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd1,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd2,2'd2,2'd1,2'd3,2'd3,2'd1,2'd1,2'd3},
'{2'd2,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_22_31[7:0][7:0] = '{'{2'd2,2'd2,2'd1,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd1,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_22_32[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2}};

parameter bit [1:0] SpriteTableB_22_33[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_22_34[7:0][7:0] = '{'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_22_35[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_23_0[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_23_1[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_23_2[7:0][7:0] = '{'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_23_3[7:0][7:0] = '{'{2'd1,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_23_4[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_23_5[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2}};

parameter bit [1:0] SpriteTableB_23_6[7:0][7:0] = '{'{2'd1,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd1},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_23_7[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_23_8[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd2,2'd2}};

parameter bit [1:0] SpriteTableB_23_9[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd1,2'd3,2'd2,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd1,2'd3,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd1,2'd3,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd2,2'd2}};

parameter bit [1:0] SpriteTableB_23_10[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd2},
'{2'd3,2'd1,2'd3,2'd3,2'd2,2'd3,2'd3,2'd2},
'{2'd3,2'd1,2'd3,2'd2,2'd2,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_23_11[7:0][7:0] = '{'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_23_12[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_23_13[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_23_14[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_23_15[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_23_16[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_23_17[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_23_18[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd2,2'd1,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd1,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_23_19[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_23_20[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_23_21[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_23_22[7:0][7:0] = '{'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_23_23[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_23_24[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_23_25[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_23_26[7:0][7:0] = '{'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd2,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_23_27[7:0][7:0] = '{'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_23_28[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd2,2'd1,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_23_29[7:0][7:0] = '{'{2'd1,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_23_30[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_23_31[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_23_32[7:0][7:0] = '{'{2'd2,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd2,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_23_33[7:0][7:0] = '{'{2'd2,2'd3,2'd3,2'd3,2'd2,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_23_34[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_23_35[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_24_0[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd2,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_24_1[7:0][7:0] = '{'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_24_2[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_24_3[7:0][7:0] = '{'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_24_4[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_24_5[7:0][7:0] = '{'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_24_6[7:0][7:0] = '{'{2'd3,2'd1,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_24_7[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd1,2'd3,2'd3,2'd3,2'd1,2'd2,2'd3,2'd3},
'{2'd3,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_24_8[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd2,2'd2,2'd3,2'd2,2'd2,2'd3,2'd2}};

parameter bit [1:0] SpriteTableB_24_9[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd2,2'd2,2'd3,2'd2,2'd2,2'd3,2'd2},
'{2'd3,2'd2,2'd2,2'd3,2'd2,2'd2,2'd3,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd3,2'd2,2'd2,2'd3}};

parameter bit [1:0] SpriteTableB_24_10[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd2,2'd2,2'd2,2'd3,2'd2,2'd2,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd2,2'd2,2'd2,2'd3},
'{2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3},
'{2'd3,2'd2,2'd2,2'd2,2'd3,2'd2,2'd2,2'd1},
'{2'd3,2'd3,2'd2,2'd2,2'd3,2'd2,2'd3,2'd1},
'{2'd3,2'd2,2'd2,2'd2,2'd3,2'd2,2'd3,2'd1},
'{2'd3,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_24_11[7:0][7:0] = '{'{2'd3,2'd3,2'd2,2'd2,2'd3,2'd2,2'd3,2'd1},
'{2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3},
'{2'd3,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd2,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_24_12[7:0][7:0] = '{'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd2,2'd3,2'd2,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_24_13[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_24_14[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_24_15[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_24_16[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_24_17[7:0][7:0] = '{'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd1,2'd1,2'd1,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_24_18[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_24_19[7:0][7:0] = '{'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_24_20[7:0][7:0] = '{'{2'd1,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_24_21[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd1,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_24_22[7:0][7:0] = '{'{2'd3,2'd2,2'd3,2'd2,2'd1,2'd1,2'd3,2'd3},
'{2'd2,2'd3,2'd2,2'd3,2'd2,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd2,2'd3,2'd1},
'{2'd3,2'd2,2'd3,2'd3,2'd2,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd2,2'd3,2'd2},
'{2'd2,2'd3,2'd2,2'd3,2'd2,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_24_23[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd2,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd2,2'd2,2'd3,2'd2,2'd3}};

parameter bit [1:0] SpriteTableB_24_24[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd1,2'd2,2'd3,2'd2,2'd1,2'd2},
'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd3},
'{2'd1,2'd3,2'd1,2'd3,2'd2,2'd2,2'd2,2'd2}};

parameter bit [1:0] SpriteTableB_24_25[7:0][7:0] = '{'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd2,2'd2},
'{2'd1,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_24_26[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_24_27[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd1,2'd2},
'{2'd3,2'd3,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd1,2'd2,2'd2,2'd2,2'd2}};

parameter bit [1:0] SpriteTableB_24_28[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd2,2'd2},
'{2'd1,2'd3,2'd3,2'd2,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd1,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_24_29[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_24_30[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_24_31[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_24_32[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_24_33[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd1,2'd3,2'd1,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_24_34[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_24_35[7:0][7:0] = '{'{2'd2,2'd3,2'd3,2'd3,2'd1,2'd1,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_25_0[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_25_1[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd1,2'd2,2'd2},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_25_2[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_25_3[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd1,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_25_4[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_25_5[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd2},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2}};

parameter bit [1:0] SpriteTableB_25_6[7:0][7:0] = '{'{2'd1,2'd3,2'd1,2'd3,2'd1,2'd3,2'd3,2'd2},
'{2'd1,2'd3,2'd1,2'd3,2'd2,2'd3,2'd3,2'd2},
'{2'd3,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd3,2'd2,2'd2,2'd2,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd3},
'{2'd1,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_25_7[7:0][7:0] = '{'{2'd2,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2}};

parameter bit [1:0] SpriteTableB_25_8[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2}};

parameter bit [1:0] SpriteTableB_25_9[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_25_10[7:0][7:0] = '{'{2'd1,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_25_11[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd2,2'd3,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd2,2'd3}};

parameter bit [1:0] SpriteTableB_25_12[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_25_13[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_25_14[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd1,2'd3,2'd1,2'd1,2'd1,2'd1},
'{2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_25_15[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_25_16[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_25_17[7:0][7:0] = '{'{2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_25_18[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_25_19[7:0][7:0] = '{'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_25_20[7:0][7:0] = '{'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_25_21[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd1,2'd3,2'd1,2'd2,2'd2,2'd3}};

parameter bit [1:0] SpriteTableB_25_22[7:0][7:0] = '{'{2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd3,2'd1},
'{2'd1,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1},
'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd1,2'd1},
'{2'd2,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd1,2'd1,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_25_23[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3},
'{2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd1,2'd1},
'{2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd1},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_25_24[7:0][7:0] = '{'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd2,2'd2,2'd2,2'd3,2'd1,2'd3,2'd1,2'd3},
'{2'd2,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd1,2'd1,2'd1,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_25_25[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd2,2'd1,2'd1,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd3,2'd3},
'{2'd3,2'd2,2'd2,2'd2,2'd3,2'd1,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd1,2'd1}};

parameter bit [1:0] SpriteTableB_25_26[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd1,2'd1,2'd1},
'{2'd1,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd1,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd1,2'd1}};

parameter bit [1:0] SpriteTableB_25_27[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_25_28[7:0][7:0] = '{'{2'd2,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_25_29[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_25_30[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_25_31[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_25_32[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_25_33[7:0][7:0] = '{'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2}};

parameter bit [1:0] SpriteTableB_25_34[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1},
'{2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd3},
'{2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd2,2'd2,2'd1,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_25_35[7:0][7:0] = '{'{2'd3,2'd3,2'd2,2'd2,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_26_0[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_26_1[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd1,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd3},
'{2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1},
'{2'd3,2'd3,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2}};

parameter bit [1:0] SpriteTableB_26_2[7:0][7:0] = '{'{2'd3,2'd2,2'd3,2'd2,2'd2,2'd2,2'd2,2'd1},
'{2'd3,2'd1,2'd1,2'd2,2'd1,2'd2,2'd1,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_26_3[7:0][7:0] = '{'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd2,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_26_4[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_26_5[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd1,2'd1,2'd1,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2}};

parameter bit [1:0] SpriteTableB_26_6[7:0][7:0] = '{'{2'd2,2'd2,2'd3,2'd1,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd2},
'{2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd2,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2}};

parameter bit [1:0] SpriteTableB_26_7[7:0][7:0] = '{'{2'd2,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd2,2'd2,2'd1,2'd1,2'd1,2'd1},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3}};

parameter bit [1:0] SpriteTableB_26_8[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd1},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd1},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_26_9[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd3,2'd2,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_26_10[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd3,2'd2,2'd2,2'd2,2'd3,2'd2,2'd2},
'{2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2}};

parameter bit [1:0] SpriteTableB_26_11[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd1,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_26_12[7:0][7:0] = '{'{2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_26_13[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_26_14[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2}};

parameter bit [1:0] SpriteTableB_26_15[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_26_16[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_26_17[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_26_18[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd2,2'd1,2'd1,2'd3,2'd2},
'{2'd3,2'd3,2'd2,2'd3,2'd2,2'd2,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_26_19[7:0][7:0] = '{'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2}};

parameter bit [1:0] SpriteTableB_26_20[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_26_21[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3}};

parameter bit [1:0] SpriteTableB_26_22[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd1,2'd3,2'd3,2'd1,2'd2},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd1,2'd3,2'd1,2'd3,2'd1,2'd1,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2},
'{2'd1,2'd1,2'd1,2'd3,2'd3,2'd1,2'd3,2'd2},
'{2'd3,2'd1,2'd1,2'd1,2'd1,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_26_23[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd1,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd1,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_26_24[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd1,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_26_25[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_26_26[7:0][7:0] = '{'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd1,2'd1,2'd1,2'd3,2'd3,2'd1,2'd1,2'd1},
'{2'd3,2'd3,2'd1,2'd1,2'd1,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd3}};

parameter bit [1:0] SpriteTableB_26_27[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1},
'{2'd3,2'd3,2'd1,2'd1,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_26_28[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_26_29[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_26_30[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_26_31[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_26_32[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_26_33[7:0][7:0] = '{'{2'd3,2'd3,2'd1,2'd2,2'd2,2'd1,2'd3,2'd3},
'{2'd3,2'd1,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3},
'{2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2}};

parameter bit [1:0] SpriteTableB_26_34[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_26_35[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_27_0[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_27_1[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_27_2[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_27_3[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd1,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd1,2'd2,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd2,2'd2,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_27_4[7:0][7:0] = '{'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_27_5[7:0][7:0] = '{'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd1,2'd1},
'{2'd1,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd1,2'd3,2'd3,2'd3,2'd1,2'd2,2'd3}};

parameter bit [1:0] SpriteTableB_27_6[7:0][7:0] = '{'{2'd2,2'd2,2'd1,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd1}};

parameter bit [1:0] SpriteTableB_27_7[7:0][7:0] = '{'{2'd1,2'd1,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_27_8[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3,2'd2}};

parameter bit [1:0] SpriteTableB_27_9[7:0][7:0] = '{'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_27_10[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd1,2'd3},
'{2'd2,2'd1,2'd1,2'd1,2'd2,2'd2,2'd1,2'd2},
'{2'd2,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd1,2'd1,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_27_11[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_27_12[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3}};

parameter bit [1:0] SpriteTableB_27_13[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd2,2'd1,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd2},
'{2'd2,2'd3,2'd3,2'd2,2'd2,2'd2,2'd3,2'd3},
'{2'd2,2'd3,2'd1,2'd2,2'd2,2'd3,2'd2,2'd3}};

parameter bit [1:0] SpriteTableB_27_14[7:0][7:0] = '{'{2'd3,2'd2,2'd3,2'd3,2'd2,2'd1,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd2,2'd2},
'{2'd2,2'd3,2'd2,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_27_15[7:0][7:0] = '{'{2'd2,2'd2,2'd3,2'd3,2'd2,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd2,2'd3,2'd3,2'd2,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_27_16[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_27_17[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd3}};

parameter bit [1:0] SpriteTableB_27_18[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd2,2'd3,2'd3,2'd2},
'{2'd2,2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd3},
'{2'd2,2'd3,2'd2,2'd2,2'd3,2'd2,2'd3,2'd2},
'{2'd2,2'd3,2'd2,2'd2,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd1,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_27_19[7:0][7:0] = '{'{2'd3,2'd2,2'd2,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd1,2'd3,2'd2,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd3,2'd3},
'{2'd3,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd2,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd1,2'd2,2'd3,2'd3,2'd2,2'd3,2'd1},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_27_20[7:0][7:0] = '{'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd2,2'd2,2'd2,2'd1},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd1,2'd1,2'd1,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_27_21[7:0][7:0] = '{'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd2,2'd2,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_27_22[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_27_23[7:0][7:0] = '{'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_27_24[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_27_25[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd1,2'd3,2'd1,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_27_26[7:0][7:0] = '{'{2'd3,2'd1,2'd3,2'd1,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd1},
'{2'd3,2'd3,2'd1,2'd2,2'd1,2'd1,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_27_27[7:0][7:0] = '{'{2'd1,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd1,2'd1,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_27_28[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_27_29[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_27_30[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_27_31[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_27_32[7:0][7:0] = '{'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd1,2'd1,2'd3,2'd3,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_27_33[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2},
'{2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_27_34[7:0][7:0] = '{'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd2,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_27_35[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_28_0[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_28_1[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1}};

parameter bit [1:0] SpriteTableB_28_2[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_28_3[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_28_4[7:0][7:0] = '{'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd2,2'd2,2'd3,2'd3,2'd1,2'd2},
'{2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1}};

parameter bit [1:0] SpriteTableB_28_5[7:0][7:0] = '{'{2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1},
'{2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1},
'{2'd3,2'd3,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd2,2'd1,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_28_6[7:0][7:0] = '{'{2'd3,2'd3,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_28_7[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd2,2'd2},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2},
'{2'd2,2'd1,2'd3,2'd3,2'd1,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd1,2'd2,2'd3,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd1,2'd1},
'{2'd3,2'd2,2'd2,2'd2,2'd2,2'd1,2'd3,2'd3},
'{2'd3,2'd2,2'd2,2'd2,2'd2,2'd1,2'd3,2'd3},
'{2'd3,2'd1,2'd2,2'd2,2'd2,2'd1,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_28_8[7:0][7:0] = '{'{2'd3,2'd1,2'd2,2'd2,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3},
'{2'd2,2'd1,2'd2,2'd1,2'd1,2'd1,2'd1,2'd1},
'{2'd2,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_28_9[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd1,2'd3,2'd3,2'd2,2'd1},
'{2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd2,2'd1,2'd3,2'd3,2'd2,2'd2,2'd3},
'{2'd3,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd2,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd1,2'd1},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd2,2'd2,2'd3,2'd3,2'd2,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_28_10[7:0][7:0] = '{'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd1,2'd3,2'd2},
'{2'd3,2'd3,2'd2,2'd2,2'd3,2'd2,2'd2,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd1,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_28_11[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd1,2'd3,2'd1,2'd3,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2}};

parameter bit [1:0] SpriteTableB_28_12[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd2,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_28_13[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd2,2'd2,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd2,2'd1,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd1,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd1,2'd1,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_28_14[7:0][7:0] = '{'{2'd2,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd1,2'd1,2'd1,2'd1,2'd3},
'{2'd3,2'd2,2'd1,2'd2,2'd3,2'd2,2'd2,2'd3},
'{2'd2,2'd2,2'd2,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd2,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_28_15[7:0][7:0] = '{'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd2},
'{2'd3,2'd2,2'd2,2'd3,2'd3,2'd2,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_28_16[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd3}};

parameter bit [1:0] SpriteTableB_28_17[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd3,2'd3},
'{2'd3,2'd2,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd1,2'd1,2'd2,2'd2,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_28_18[7:0][7:0] = '{'{2'd3,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd2,2'd1,2'd3,2'd1,2'd2,2'd3,2'd3,2'd1},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd3,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2}};

parameter bit [1:0] SpriteTableB_28_19[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd2},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_28_20[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd1,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd3,2'd1,2'd3,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd2,2'd2,2'd3,2'd2,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_28_21[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd2,2'd3,2'd3},
'{2'd2,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd2,2'd2,2'd3,2'd3,2'd2,2'd2}};

parameter bit [1:0] SpriteTableB_28_22[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_28_23[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1}};

parameter bit [1:0] SpriteTableB_28_24[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_28_25[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd1,2'd2},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd2,2'd1,2'd1},
'{2'd1,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd1},
'{2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2}};

parameter bit [1:0] SpriteTableB_28_26[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd1,2'd1,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_28_27[7:0][7:0] = '{'{2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_28_28[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_28_29[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_28_30[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_28_31[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_28_32[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_28_33[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_28_34[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd2,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_28_35[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_29_0[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_29_1[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_29_2[7:0][7:0] = '{'{2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_29_3[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_29_4[7:0][7:0] = '{'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd1,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_29_5[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_29_6[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd1,2'd2,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd2,2'd2,2'd1,2'd3},
'{2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd1},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd1,2'd1}};

parameter bit [1:0] SpriteTableB_29_7[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd2,2'd3,2'd3,2'd2,2'd1,2'd2,2'd2,2'd2},
'{2'd1,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_29_8[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_29_9[7:0][7:0] = '{'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1},
'{2'd3,2'd3,2'd2,2'd3,2'd2,2'd2,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_29_10[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd3,2'd3,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3,2'd2},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd2,2'd2,2'd3,2'd2,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd2,2'd3,2'd2}};

parameter bit [1:0] SpriteTableB_29_11[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd2,2'd3,2'd2,2'd3,2'd2,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd3,2'd2,2'd2,2'd2,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_29_12[7:0][7:0] = '{'{2'd3,2'd3,2'd1,2'd2,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd2,2'd3,2'd3,2'd1,2'd3,2'd1,2'd3,2'd2},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_29_13[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd2},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_29_14[7:0][7:0] = '{'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2}};

parameter bit [1:0] SpriteTableB_29_15[7:0][7:0] = '{'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd2,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd1,2'd1,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_29_16[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2},
'{2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_29_17[7:0][7:0] = '{'{2'd3,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd3,2'd3},
'{2'd3,2'd2,2'd2,2'd3,2'd2,2'd2,2'd2,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd2,2'd2,2'd1,2'd3,2'd3,2'd1},
'{2'd3,2'd1,2'd2,2'd1,2'd1,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_29_18[7:0][7:0] = '{'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_29_19[7:0][7:0] = '{'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd1,2'd3,2'd3,2'd3,2'd1,2'd1}};

parameter bit [1:0] SpriteTableB_29_20[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd1,2'd1,2'd2,2'd2,2'd1},
'{2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3},
'{2'd3,2'd1,2'd2,2'd2,2'd2,2'd2,2'd1,2'd3},
'{2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd1,2'd3},
'{2'd1,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3},
'{2'd2,2'd1,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2}};

parameter bit [1:0] SpriteTableB_29_21[7:0][7:0] = '{'{2'd3,2'd2,2'd2,2'd2,2'd3,2'd1,2'd3,2'd3},
'{2'd3,2'd2,2'd2,2'd3,2'd2,2'd1,2'd3,2'd3},
'{2'd3,2'd2,2'd2,2'd3,2'd3,2'd1,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd1},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd1,2'd2},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2},
'{2'd2,2'd3,2'd3,2'd2,2'd3,2'd3,2'd2,2'd2}};

parameter bit [1:0] SpriteTableB_29_22[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd3,2'd2},
'{2'd2,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd2,2'd1}};

parameter bit [1:0] SpriteTableB_29_23[7:0][7:0] = '{'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd1,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd2,2'd1,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd2,2'd2,2'd2},
'{2'd1,2'd1,2'd2,2'd1,2'd3,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_29_24[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3},
'{2'd1,2'd1,2'd3,2'd2,2'd3,2'd3,2'd3,2'd1},
'{2'd1,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_29_25[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3,2'd2},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_29_26[7:0][7:0] = '{'{2'd2,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1}};

parameter bit [1:0] SpriteTableB_29_27[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_29_28[7:0][7:0] = '{'{2'd3,2'd3,2'd2,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd2,2'd2,2'd2,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_29_29[7:0][7:0] = '{'{2'd3,2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_29_30[7:0][7:0] = '{'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_29_31[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_29_32[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_29_33[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_29_34[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_29_35[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_30_0[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_30_1[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd1,2'd1,2'd3},
'{2'd3,2'd3,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1},
'{2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_30_2[7:0][7:0] = '{'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_30_3[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_30_4[7:0][7:0] = '{'{2'd1,2'd3,2'd1,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd1,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_30_5[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_30_6[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_30_7[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_30_8[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd1,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_30_9[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd1,2'd2,2'd2},
'{2'd3,2'd3,2'd1,2'd2,2'd2,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2,2'd3}};

parameter bit [1:0] SpriteTableB_30_10[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd1,2'd2,2'd1,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd2,2'd1,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_30_11[7:0][7:0] = '{'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd2},
'{2'd2,2'd2,2'd2,2'd1,2'd2,2'd3,2'd3,2'd2},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd1,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_30_12[7:0][7:0] = '{'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd2,2'd2,2'd3,2'd1,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_30_13[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd1,2'd2},
'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd1,2'd2}};

parameter bit [1:0] SpriteTableB_30_14[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_30_15[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd2},
'{2'd2,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd1,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd1,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_30_16[7:0][7:0] = '{'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd1,2'd3},
'{2'd2,2'd3,2'd3,2'd2,2'd2,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd2,2'd3,2'd3,2'd3,2'd2,2'd2,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_30_17[7:0][7:0] = '{'{2'd3,2'd3,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd1,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd2,2'd2,2'd2,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd2,2'd3,2'd3},
'{2'd2,2'd3,2'd1,2'd3,2'd2,2'd3,2'd1,2'd3},
'{2'd1,2'd2,2'd1,2'd3,2'd1,2'd3,2'd2,2'd3}};

parameter bit [1:0] SpriteTableB_30_18[7:0][7:0] = '{'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3}};

parameter bit [1:0] SpriteTableB_30_19[7:0][7:0] = '{'{2'd3,2'd3,2'd1,2'd1,2'd1,2'd1,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd1},
'{2'd3,2'd3,2'd3,2'd1,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd1,2'd2,2'd2,2'd2,2'd2},
'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd2,2'd2,2'd1},
'{2'd3,2'd3,2'd1,2'd1,2'd1,2'd1,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_30_20[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_30_21[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_30_22[7:0][7:0] = '{'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd2,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd1,2'd2,2'd3,2'd2,2'd1,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_30_23[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_30_24[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_30_25[7:0][7:0] = '{'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_30_26[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_30_27[7:0][7:0] = '{'{2'd3,2'd3,2'd2,2'd2,2'd1,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_30_28[7:0][7:0] = '{'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_30_29[7:0][7:0] = '{'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_30_30[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_30_31[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_30_32[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_30_33[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_30_34[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_30_35[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_31_0[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_31_1[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_31_2[7:0][7:0] = '{'{2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_31_3[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_31_4[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_31_5[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_31_6[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_31_7[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_31_8[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_31_9[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd1},
'{2'd3,2'd3,2'd3,2'd3,2'd1,2'd2,2'd2,2'd3},
'{2'd3,2'd1,2'd2,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_31_10[7:0][7:0] = '{'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_31_11[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd1,2'd1,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_31_12[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd2,2'd3,2'd2,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd2,2'd3,2'd3},
'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd1,2'd3},
'{2'd3,2'd1,2'd3,2'd2,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_31_13[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd2,2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_31_14[7:0][7:0] = '{'{2'd2,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_31_15[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_31_16[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd2,2'd2,2'd1,2'd3,2'd3},
'{2'd3,2'd3,2'd2,2'd2,2'd1,2'd3,2'd3,2'd3},
'{2'd2,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_31_17[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_31_18[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_31_19[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_31_20[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_31_21[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_31_22[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_31_23[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_31_24[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_31_25[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_31_26[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_31_27[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd1,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_31_28[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_31_29[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_31_30[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_31_31[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_31_32[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_31_33[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_31_34[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

parameter bit [1:0] SpriteTableB_31_35[7:0][7:0] = '{'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3},
'{2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3,2'd3}};

assign SpriteR = SpritePaletteR[SpriteTableR];
assign SpriteG = SpritePaletteG[SpriteTableG];
assign SpriteB = SpritePaletteB[SpriteTableB];

endmodule
