//module scoreboard (
//	input logic Clk,
//	input logic Reset,
//);
//
//endmodule
