module cookies_wrapper_all (
	input logic Reset,
	input logic Clk,
	input logic [9:0] BallX,
	input logic [9:0] BallY,
	input logic [9:0] Ball_Size,

	output logic [240:0] Not_ate
);

cookie ck0 (.Clk(Clk), .Reset(Reset), .Xc(10'd498), .Yc(10'd428), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[0]) );

cookie ck1 (.Clk(Clk), .Reset(Reset), .Xc(10'd483), .Yc(10'd428), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[1]) );

cookie ck2 (.Clk(Clk), .Reset(Reset), .Xc(10'd469), .Yc(10'd428), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[2]) );

cookie ck3 (.Clk(Clk), .Reset(Reset), .Xc(10'd455), .Yc(10'd428), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[3]) );

cookie ck4 (.Clk(Clk), .Reset(Reset), .Xc(10'd441), .Yc(10'd428), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[4]) );

cookie ck5 (.Clk(Clk), .Reset(Reset), .Xc(10'd426), .Yc(10'd428), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[5]) );

cookie ck6 (.Clk(Clk), .Reset(Reset), .Xc(10'd412), .Yc(10'd428), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[6]) );

cookie ck7 (.Clk(Clk), .Reset(Reset), .Xc(10'd398), .Yc(10'd428), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[7]) );

cookie ck8 (.Clk(Clk), .Reset(Reset), .Xc(10'd383), .Yc(10'd428), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[8]) );

cookie ck9 (.Clk(Clk), .Reset(Reset), .Xc(10'd369), .Yc(10'd428), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[9]) );

cookie ck10 (.Clk(Clk), .Reset(Reset), .Xc(10'd355), .Yc(10'd428), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[10]) );

cookie ck11 (.Clk(Clk), .Reset(Reset), .Xc(10'd341), .Yc(10'd428), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[11]) );

cookie ck12 (.Clk(Clk), .Reset(Reset), .Xc(10'd326), .Yc(10'd428), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[12]) );

cookie ck13 (.Clk(Clk), .Reset(Reset), .Xc(10'd312), .Yc(10'd428), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[13]) );

cookie ck14 (.Clk(Clk), .Reset(Reset), .Xc(10'd298), .Yc(10'd428), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[14]) );

cookie ck15 (.Clk(Clk), .Reset(Reset), .Xc(10'd283), .Yc(10'd428), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[15]) );

cookie ck16 (.Clk(Clk), .Reset(Reset), .Xc(10'd269), .Yc(10'd428), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[16]) );

cookie ck17 (.Clk(Clk), .Reset(Reset), .Xc(10'd255), .Yc(10'd428), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[17]) );

cookie ck18 (.Clk(Clk), .Reset(Reset), .Xc(10'd241), .Yc(10'd428), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[18]) );

cookie ck19 (.Clk(Clk), .Reset(Reset), .Xc(10'd226), .Yc(10'd428), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[19]) );

cookie ck20 (.Clk(Clk), .Reset(Reset), .Xc(10'd212), .Yc(10'd428), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[20]) );

cookie ck21 (.Clk(Clk), .Reset(Reset), .Xc(10'd198), .Yc(10'd428), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[21]) );

cookie ck22 (.Clk(Clk), .Reset(Reset), .Xc(10'd183), .Yc(10'd428), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[22]) );

cookie ck23 (.Clk(Clk), .Reset(Reset), .Xc(10'd169), .Yc(10'd428), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[23]) );

cookie ck24 (.Clk(Clk), .Reset(Reset), .Xc(10'd155), .Yc(10'd428), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[24]) );

cookie ck25 (.Clk(Clk), .Reset(Reset), .Xc(10'd141), .Yc(10'd428), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[25]) );

cookie ck26 (.Clk(Clk), .Reset(Reset), .Xc(10'd498), .Yc(10'd415), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[26]) );

cookie ck27 (.Clk(Clk), .Reset(Reset), .Xc(10'd341), .Yc(10'd415), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[27]) );

cookie ck28 (.Clk(Clk), .Reset(Reset), .Xc(10'd298), .Yc(10'd415), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[28]) );

cookie ck29 (.Clk(Clk), .Reset(Reset), .Xc(10'd141), .Yc(10'd415), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[29]) );

cookie ck30 (.Clk(Clk), .Reset(Reset), .Xc(10'd498), .Yc(10'd402), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[30]) );

cookie ck31 (.Clk(Clk), .Reset(Reset), .Xc(10'd341), .Yc(10'd402), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[31]) );

cookie ck32 (.Clk(Clk), .Reset(Reset), .Xc(10'd298), .Yc(10'd402), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[32]) );

cookie ck33 (.Clk(Clk), .Reset(Reset), .Xc(10'd141), .Yc(10'd402), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[33]) );

cookie ck34 (.Clk(Clk), .Reset(Reset), .Xc(10'd498), .Yc(10'd389), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[34]) );

cookie ck35 (.Clk(Clk), .Reset(Reset), .Xc(10'd483), .Yc(10'd389), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[35]) );

cookie ck36 (.Clk(Clk), .Reset(Reset), .Xc(10'd469), .Yc(10'd389), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[36]) );

cookie ck37 (.Clk(Clk), .Reset(Reset), .Xc(10'd455), .Yc(10'd389), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[37]) );

cookie ck38 (.Clk(Clk), .Reset(Reset), .Xc(10'd441), .Yc(10'd389), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[38]) );

cookie ck39 (.Clk(Clk), .Reset(Reset), .Xc(10'd426), .Yc(10'd389), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[39]) );

cookie ck40 (.Clk(Clk), .Reset(Reset), .Xc(10'd383), .Yc(10'd389), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[40]) );

cookie ck41 (.Clk(Clk), .Reset(Reset), .Xc(10'd369), .Yc(10'd389), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[41]) );

cookie ck42 (.Clk(Clk), .Reset(Reset), .Xc(10'd355), .Yc(10'd389), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[42]) );

cookie ck43 (.Clk(Clk), .Reset(Reset), .Xc(10'd341), .Yc(10'd389), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[43]) );

cookie ck44 (.Clk(Clk), .Reset(Reset), .Xc(10'd298), .Yc(10'd389), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[44]) );

cookie ck45 (.Clk(Clk), .Reset(Reset), .Xc(10'd283), .Yc(10'd389), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[45]) );

cookie ck46 (.Clk(Clk), .Reset(Reset), .Xc(10'd269), .Yc(10'd389), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[46]) );

cookie ck47 (.Clk(Clk), .Reset(Reset), .Xc(10'd255), .Yc(10'd389), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[47]) );

cookie ck48 (.Clk(Clk), .Reset(Reset), .Xc(10'd212), .Yc(10'd389), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[48]) );

cookie ck49 (.Clk(Clk), .Reset(Reset), .Xc(10'd198), .Yc(10'd389), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[49]) );

cookie ck50 (.Clk(Clk), .Reset(Reset), .Xc(10'd183), .Yc(10'd389), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[50]) );

cookie ck51 (.Clk(Clk), .Reset(Reset), .Xc(10'd169), .Yc(10'd389), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[51]) );

cookie ck52 (.Clk(Clk), .Reset(Reset), .Xc(10'd155), .Yc(10'd389), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[52]) );

cookie ck53 (.Clk(Clk), .Reset(Reset), .Xc(10'd141), .Yc(10'd389), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[53]) );

cookie ck54 (.Clk(Clk), .Reset(Reset), .Xc(10'd469), .Yc(10'd376), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[54]) );

cookie ck55 (.Clk(Clk), .Reset(Reset), .Xc(10'd426), .Yc(10'd376), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[55]) );

cookie ck56 (.Clk(Clk), .Reset(Reset), .Xc(10'd383), .Yc(10'd376), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[56]) );

cookie ck57 (.Clk(Clk), .Reset(Reset), .Xc(10'd255), .Yc(10'd376), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[57]) );

cookie ck58 (.Clk(Clk), .Reset(Reset), .Xc(10'd212), .Yc(10'd376), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[58]) );

cookie ck59 (.Clk(Clk), .Reset(Reset), .Xc(10'd169), .Yc(10'd376), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[59]) );

cookie ck60 (.Clk(Clk), .Reset(Reset), .Xc(10'd469), .Yc(10'd364), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[60]) );

cookie ck61 (.Clk(Clk), .Reset(Reset), .Xc(10'd426), .Yc(10'd364), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[61]) );

cookie ck62 (.Clk(Clk), .Reset(Reset), .Xc(10'd383), .Yc(10'd364), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[62]) );

cookie ck63 (.Clk(Clk), .Reset(Reset), .Xc(10'd255), .Yc(10'd364), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[63]) );

cookie ck64 (.Clk(Clk), .Reset(Reset), .Xc(10'd212), .Yc(10'd364), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[64]) );

cookie ck65 (.Clk(Clk), .Reset(Reset), .Xc(10'd169), .Yc(10'd364), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[65]) );

cookie ck66 (.Clk(Clk), .Reset(Reset), .Xc(10'd483), .Yc(10'd351), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[66]) );

cookie ck67 (.Clk(Clk), .Reset(Reset), .Xc(10'd469), .Yc(10'd351), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[67]) );

cookie ck68 (.Clk(Clk), .Reset(Reset), .Xc(10'd426), .Yc(10'd351), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[68]) );

cookie ck69 (.Clk(Clk), .Reset(Reset), .Xc(10'd412), .Yc(10'd351), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[69]) );

cookie ck70 (.Clk(Clk), .Reset(Reset), .Xc(10'd398), .Yc(10'd351), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[70]) );

cookie ck71 (.Clk(Clk), .Reset(Reset), .Xc(10'd383), .Yc(10'd351), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[71]) );

cookie ck72 (.Clk(Clk), .Reset(Reset), .Xc(10'd369), .Yc(10'd351), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[72]) );

cookie ck73 (.Clk(Clk), .Reset(Reset), .Xc(10'd355), .Yc(10'd351), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[73]) );

cookie ck74 (.Clk(Clk), .Reset(Reset), .Xc(10'd341), .Yc(10'd351), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[74]) );

cookie ck75 (.Clk(Clk), .Reset(Reset), .Xc(10'd298), .Yc(10'd351), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[75]) );

cookie ck76 (.Clk(Clk), .Reset(Reset), .Xc(10'd283), .Yc(10'd351), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[76]) );

cookie ck77 (.Clk(Clk), .Reset(Reset), .Xc(10'd269), .Yc(10'd351), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[77]) );

cookie ck78 (.Clk(Clk), .Reset(Reset), .Xc(10'd255), .Yc(10'd351), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[78]) );

cookie ck79 (.Clk(Clk), .Reset(Reset), .Xc(10'd241), .Yc(10'd351), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[79]) );

cookie ck80 (.Clk(Clk), .Reset(Reset), .Xc(10'd226), .Yc(10'd351), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[80]) );

cookie ck81 (.Clk(Clk), .Reset(Reset), .Xc(10'd212), .Yc(10'd351), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[81]) );

cookie ck82 (.Clk(Clk), .Reset(Reset), .Xc(10'd169), .Yc(10'd351), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[82]) );

cookie ck83 (.Clk(Clk), .Reset(Reset), .Xc(10'd155), .Yc(10'd351), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[83]) );

cookie ck84 (.Clk(Clk), .Reset(Reset), .Xc(10'd498), .Yc(10'd338), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[84]) );

cookie ck85 (.Clk(Clk), .Reset(Reset), .Xc(10'd426), .Yc(10'd338), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[85]) );

cookie ck86 (.Clk(Clk), .Reset(Reset), .Xc(10'd341), .Yc(10'd338), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[86]) );

cookie ck87 (.Clk(Clk), .Reset(Reset), .Xc(10'd298), .Yc(10'd338), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[87]) );

cookie ck88 (.Clk(Clk), .Reset(Reset), .Xc(10'd212), .Yc(10'd338), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[88]) );

cookie ck89 (.Clk(Clk), .Reset(Reset), .Xc(10'd141), .Yc(10'd338), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[89]) );

cookie ck90 (.Clk(Clk), .Reset(Reset), .Xc(10'd498), .Yc(10'd325), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[90]) );

cookie ck91 (.Clk(Clk), .Reset(Reset), .Xc(10'd426), .Yc(10'd325), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[91]) );

cookie ck92 (.Clk(Clk), .Reset(Reset), .Xc(10'd341), .Yc(10'd325), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[92]) );

cookie ck93 (.Clk(Clk), .Reset(Reset), .Xc(10'd298), .Yc(10'd325), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[93]) );

cookie ck94 (.Clk(Clk), .Reset(Reset), .Xc(10'd212), .Yc(10'd325), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[94]) );

cookie ck95 (.Clk(Clk), .Reset(Reset), .Xc(10'd141), .Yc(10'd325), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[95]) );

cookie ck96 (.Clk(Clk), .Reset(Reset), .Xc(10'd498), .Yc(10'd312), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[96]) );

cookie ck97 (.Clk(Clk), .Reset(Reset), .Xc(10'd483), .Yc(10'd312), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[97]) );

cookie ck98 (.Clk(Clk), .Reset(Reset), .Xc(10'd469), .Yc(10'd312), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[98]) );

cookie ck99 (.Clk(Clk), .Reset(Reset), .Xc(10'd455), .Yc(10'd312), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[99]) );

cookie ck100 (.Clk(Clk), .Reset(Reset), .Xc(10'd441), .Yc(10'd312), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[100]) );

cookie ck101 (.Clk(Clk), .Reset(Reset), .Xc(10'd426), .Yc(10'd312), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[101]) );

cookie ck102 (.Clk(Clk), .Reset(Reset), .Xc(10'd412), .Yc(10'd312), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[102]) );

cookie ck103 (.Clk(Clk), .Reset(Reset), .Xc(10'd398), .Yc(10'd312), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[103]) );

cookie ck104 (.Clk(Clk), .Reset(Reset), .Xc(10'd383), .Yc(10'd312), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[104]) );

cookie ck105 (.Clk(Clk), .Reset(Reset), .Xc(10'd369), .Yc(10'd312), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[105]) );

cookie ck106 (.Clk(Clk), .Reset(Reset), .Xc(10'd355), .Yc(10'd312), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[106]) );

cookie ck107 (.Clk(Clk), .Reset(Reset), .Xc(10'd341), .Yc(10'd312), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[107]) );

cookie ck108 (.Clk(Clk), .Reset(Reset), .Xc(10'd298), .Yc(10'd312), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[108]) );

cookie ck109 (.Clk(Clk), .Reset(Reset), .Xc(10'd283), .Yc(10'd312), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[109]) );

cookie ck110 (.Clk(Clk), .Reset(Reset), .Xc(10'd269), .Yc(10'd312), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[110]) );

cookie ck111 (.Clk(Clk), .Reset(Reset), .Xc(10'd255), .Yc(10'd312), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[111]) );

cookie ck112 (.Clk(Clk), .Reset(Reset), .Xc(10'd241), .Yc(10'd312), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[112]) );

cookie ck113 (.Clk(Clk), .Reset(Reset), .Xc(10'd226), .Yc(10'd312), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[113]) );

cookie ck114 (.Clk(Clk), .Reset(Reset), .Xc(10'd212), .Yc(10'd312), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[114]) );

cookie ck115 (.Clk(Clk), .Reset(Reset), .Xc(10'd198), .Yc(10'd312), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[115]) );

cookie ck116 (.Clk(Clk), .Reset(Reset), .Xc(10'd183), .Yc(10'd312), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[116]) );

cookie ck117 (.Clk(Clk), .Reset(Reset), .Xc(10'd169), .Yc(10'd312), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[117]) );

cookie ck118 (.Clk(Clk), .Reset(Reset), .Xc(10'd155), .Yc(10'd312), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[118]) );

cookie ck119 (.Clk(Clk), .Reset(Reset), .Xc(10'd141), .Yc(10'd312), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[119]) );

cookie ck120 (.Clk(Clk), .Reset(Reset), .Xc(10'd426), .Yc(10'd299), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[120]) );

cookie ck121 (.Clk(Clk), .Reset(Reset), .Xc(10'd212), .Yc(10'd299), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[121]) );

cookie ck122 (.Clk(Clk), .Reset(Reset), .Xc(10'd426), .Yc(10'd286), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[122]) );

cookie ck123 (.Clk(Clk), .Reset(Reset), .Xc(10'd212), .Yc(10'd286), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[123]) );

cookie ck124 (.Clk(Clk), .Reset(Reset), .Xc(10'd426), .Yc(10'd273), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[124]) );

cookie ck125 (.Clk(Clk), .Reset(Reset), .Xc(10'd212), .Yc(10'd273), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[125]) );

cookie ck126 (.Clk(Clk), .Reset(Reset), .Xc(10'd426), .Yc(10'd260), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[126]) );

cookie ck127 (.Clk(Clk), .Reset(Reset), .Xc(10'd212), .Yc(10'd260), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[127]) );

cookie ck128 (.Clk(Clk), .Reset(Reset), .Xc(10'd426), .Yc(10'd247), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[128]) );

cookie ck129 (.Clk(Clk), .Reset(Reset), .Xc(10'd212), .Yc(10'd247), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[129]) );

cookie ck130 (.Clk(Clk), .Reset(Reset), .Xc(10'd426), .Yc(10'd234), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[130]) );

cookie ck131 (.Clk(Clk), .Reset(Reset), .Xc(10'd212), .Yc(10'd234), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[131]) );

cookie ck132 (.Clk(Clk), .Reset(Reset), .Xc(10'd426), .Yc(10'd222), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[132]) );

cookie ck133 (.Clk(Clk), .Reset(Reset), .Xc(10'd212), .Yc(10'd222), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[133]) );

cookie ck134 (.Clk(Clk), .Reset(Reset), .Xc(10'd426), .Yc(10'd209), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[134]) );

cookie ck135 (.Clk(Clk), .Reset(Reset), .Xc(10'd212), .Yc(10'd209), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[135]) );

cookie ck136 (.Clk(Clk), .Reset(Reset), .Xc(10'd426), .Yc(10'd196), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[136]) );

cookie ck137 (.Clk(Clk), .Reset(Reset), .Xc(10'd212), .Yc(10'd196), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[137]) );

cookie ck138 (.Clk(Clk), .Reset(Reset), .Xc(10'd426), .Yc(10'd183), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[138]) );

cookie ck139 (.Clk(Clk), .Reset(Reset), .Xc(10'd212), .Yc(10'd183), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[139]) );

cookie ck140 (.Clk(Clk), .Reset(Reset), .Xc(10'd426), .Yc(10'd170), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[140]) );

cookie ck141 (.Clk(Clk), .Reset(Reset), .Xc(10'd212), .Yc(10'd170), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[141]) );

cookie ck142 (.Clk(Clk), .Reset(Reset), .Xc(10'd498), .Yc(10'd157), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[142]) );

cookie ck143 (.Clk(Clk), .Reset(Reset), .Xc(10'd483), .Yc(10'd157), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[143]) );

cookie ck144 (.Clk(Clk), .Reset(Reset), .Xc(10'd469), .Yc(10'd157), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[144]) );

cookie ck145 (.Clk(Clk), .Reset(Reset), .Xc(10'd455), .Yc(10'd157), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[145]) );

cookie ck146 (.Clk(Clk), .Reset(Reset), .Xc(10'd441), .Yc(10'd157), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[146]) );

cookie ck147 (.Clk(Clk), .Reset(Reset), .Xc(10'd426), .Yc(10'd157), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[147]) );

cookie ck148 (.Clk(Clk), .Reset(Reset), .Xc(10'd383), .Yc(10'd157), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[148]) );

cookie ck149 (.Clk(Clk), .Reset(Reset), .Xc(10'd369), .Yc(10'd157), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[149]) );

cookie ck150 (.Clk(Clk), .Reset(Reset), .Xc(10'd355), .Yc(10'd157), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[150]) );

cookie ck151 (.Clk(Clk), .Reset(Reset), .Xc(10'd341), .Yc(10'd157), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[151]) );

cookie ck152 (.Clk(Clk), .Reset(Reset), .Xc(10'd298), .Yc(10'd157), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[152]) );

cookie ck153 (.Clk(Clk), .Reset(Reset), .Xc(10'd283), .Yc(10'd157), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[153]) );

cookie ck154 (.Clk(Clk), .Reset(Reset), .Xc(10'd269), .Yc(10'd157), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[154]) );

cookie ck155 (.Clk(Clk), .Reset(Reset), .Xc(10'd255), .Yc(10'd157), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[155]) );

cookie ck156 (.Clk(Clk), .Reset(Reset), .Xc(10'd212), .Yc(10'd157), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[156]) );

cookie ck157 (.Clk(Clk), .Reset(Reset), .Xc(10'd198), .Yc(10'd157), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[157]) );

cookie ck158 (.Clk(Clk), .Reset(Reset), .Xc(10'd183), .Yc(10'd157), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[158]) );

cookie ck159 (.Clk(Clk), .Reset(Reset), .Xc(10'd169), .Yc(10'd157), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[159]) );

cookie ck160 (.Clk(Clk), .Reset(Reset), .Xc(10'd155), .Yc(10'd157), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[160]) );

cookie ck161 (.Clk(Clk), .Reset(Reset), .Xc(10'd141), .Yc(10'd157), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[161]) );

cookie ck162 (.Clk(Clk), .Reset(Reset), .Xc(10'd498), .Yc(10'd144), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[162]) );

cookie ck163 (.Clk(Clk), .Reset(Reset), .Xc(10'd426), .Yc(10'd144), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[163]) );

cookie ck164 (.Clk(Clk), .Reset(Reset), .Xc(10'd383), .Yc(10'd144), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[164]) );

cookie ck165 (.Clk(Clk), .Reset(Reset), .Xc(10'd255), .Yc(10'd144), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[165]) );

cookie ck166 (.Clk(Clk), .Reset(Reset), .Xc(10'd212), .Yc(10'd144), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[166]) );

cookie ck167 (.Clk(Clk), .Reset(Reset), .Xc(10'd141), .Yc(10'd144), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[167]) );

cookie ck168 (.Clk(Clk), .Reset(Reset), .Xc(10'd498), .Yc(10'd131), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[168]) );

cookie ck169 (.Clk(Clk), .Reset(Reset), .Xc(10'd426), .Yc(10'd131), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[169]) );

cookie ck170 (.Clk(Clk), .Reset(Reset), .Xc(10'd383), .Yc(10'd131), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[170]) );

cookie ck171 (.Clk(Clk), .Reset(Reset), .Xc(10'd255), .Yc(10'd131), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[171]) );

cookie ck172 (.Clk(Clk), .Reset(Reset), .Xc(10'd212), .Yc(10'd131), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[172]) );

cookie ck173 (.Clk(Clk), .Reset(Reset), .Xc(10'd141), .Yc(10'd131), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[173]) );

cookie ck174 (.Clk(Clk), .Reset(Reset), .Xc(10'd498), .Yc(10'd118), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[174]) );

cookie ck175 (.Clk(Clk), .Reset(Reset), .Xc(10'd483), .Yc(10'd118), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[175]) );

cookie ck176 (.Clk(Clk), .Reset(Reset), .Xc(10'd469), .Yc(10'd118), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[176]) );

cookie ck177 (.Clk(Clk), .Reset(Reset), .Xc(10'd455), .Yc(10'd118), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[177]) );

cookie ck178 (.Clk(Clk), .Reset(Reset), .Xc(10'd441), .Yc(10'd118), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[178]) );

cookie ck179 (.Clk(Clk), .Reset(Reset), .Xc(10'd426), .Yc(10'd118), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[179]) );

cookie ck180 (.Clk(Clk), .Reset(Reset), .Xc(10'd412), .Yc(10'd118), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[180]) );

cookie ck181 (.Clk(Clk), .Reset(Reset), .Xc(10'd398), .Yc(10'd118), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[181]) );

cookie ck182 (.Clk(Clk), .Reset(Reset), .Xc(10'd383), .Yc(10'd118), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[182]) );

cookie ck183 (.Clk(Clk), .Reset(Reset), .Xc(10'd369), .Yc(10'd118), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[183]) );

cookie ck184 (.Clk(Clk), .Reset(Reset), .Xc(10'd355), .Yc(10'd118), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[184]) );

cookie ck185 (.Clk(Clk), .Reset(Reset), .Xc(10'd341), .Yc(10'd118), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[185]) );

cookie ck186 (.Clk(Clk), .Reset(Reset), .Xc(10'd326), .Yc(10'd118), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[186]) );

cookie ck187 (.Clk(Clk), .Reset(Reset), .Xc(10'd312), .Yc(10'd118), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[187]) );

cookie ck188 (.Clk(Clk), .Reset(Reset), .Xc(10'd298), .Yc(10'd118), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[188]) );

cookie ck189 (.Clk(Clk), .Reset(Reset), .Xc(10'd283), .Yc(10'd118), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[189]) );

cookie ck190 (.Clk(Clk), .Reset(Reset), .Xc(10'd269), .Yc(10'd118), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[190]) );

cookie ck191 (.Clk(Clk), .Reset(Reset), .Xc(10'd255), .Yc(10'd118), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[191]) );

cookie ck192 (.Clk(Clk), .Reset(Reset), .Xc(10'd241), .Yc(10'd118), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[192]) );

cookie ck193 (.Clk(Clk), .Reset(Reset), .Xc(10'd226), .Yc(10'd118), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[193]) );

cookie ck194 (.Clk(Clk), .Reset(Reset), .Xc(10'd212), .Yc(10'd118), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[194]) );

cookie ck195 (.Clk(Clk), .Reset(Reset), .Xc(10'd198), .Yc(10'd118), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[195]) );

cookie ck196 (.Clk(Clk), .Reset(Reset), .Xc(10'd183), .Yc(10'd118), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[196]) );

cookie ck197 (.Clk(Clk), .Reset(Reset), .Xc(10'd169), .Yc(10'd118), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[197]) );

cookie ck198 (.Clk(Clk), .Reset(Reset), .Xc(10'd155), .Yc(10'd118), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[198]) );

cookie ck199 (.Clk(Clk), .Reset(Reset), .Xc(10'd141), .Yc(10'd118), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[199]) );

cookie ck200 (.Clk(Clk), .Reset(Reset), .Xc(10'd498), .Yc(10'd105), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[200]) );

cookie ck201 (.Clk(Clk), .Reset(Reset), .Xc(10'd341), .Yc(10'd105), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[201]) );

cookie ck202 (.Clk(Clk), .Reset(Reset), .Xc(10'd298), .Yc(10'd105), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[202]) );

cookie ck203 (.Clk(Clk), .Reset(Reset), .Xc(10'd141), .Yc(10'd105), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[203]) );

cookie ck204 (.Clk(Clk), .Reset(Reset), .Xc(10'd426), .Yc(10'd105), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[204]) );

cookie ck205 (.Clk(Clk), .Reset(Reset), .Xc(10'd212), .Yc(10'd105), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[205]) );

cookie ck206 (.Clk(Clk), .Reset(Reset), .Xc(10'd426), .Yc(10'd93), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[206]) );

cookie ck207 (.Clk(Clk), .Reset(Reset), .Xc(10'd341), .Yc(10'd93), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[207]) );

cookie ck208 (.Clk(Clk), .Reset(Reset), .Xc(10'd298), .Yc(10'd93), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[208]) );

cookie ck209 (.Clk(Clk), .Reset(Reset), .Xc(10'd212), .Yc(10'd93), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[209]) );

cookie ck210 (.Clk(Clk), .Reset(Reset), .Xc(10'd498), .Yc(10'd80), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[210]) );

cookie ck211 (.Clk(Clk), .Reset(Reset), .Xc(10'd426), .Yc(10'd80), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[211]) );

cookie ck212 (.Clk(Clk), .Reset(Reset), .Xc(10'd341), .Yc(10'd80), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[212]) );

cookie ck213 (.Clk(Clk), .Reset(Reset), .Xc(10'd298), .Yc(10'd80), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[213]) );

cookie ck214 (.Clk(Clk), .Reset(Reset), .Xc(10'd212), .Yc(10'd80), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[214]) );

cookie ck215 (.Clk(Clk), .Reset(Reset), .Xc(10'd141), .Yc(10'd80), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[215]) );

cookie ck216 (.Clk(Clk), .Reset(Reset), .Xc(10'd498), .Yc(10'd67), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[216]) );

cookie ck217 (.Clk(Clk), .Reset(Reset), .Xc(10'd483), .Yc(10'd67), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[217]) );

cookie ck218 (.Clk(Clk), .Reset(Reset), .Xc(10'd469), .Yc(10'd67), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[218]) );

cookie ck219 (.Clk(Clk), .Reset(Reset), .Xc(10'd455), .Yc(10'd67), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[219]) );

cookie ck220 (.Clk(Clk), .Reset(Reset), .Xc(10'd441), .Yc(10'd67), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[220]) );

cookie ck221 (.Clk(Clk), .Reset(Reset), .Xc(10'd426), .Yc(10'd67), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[221]) );

cookie ck222 (.Clk(Clk), .Reset(Reset), .Xc(10'd412), .Yc(10'd67), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[222]) );

cookie ck223 (.Clk(Clk), .Reset(Reset), .Xc(10'd398), .Yc(10'd67), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[223]) );

cookie ck224 (.Clk(Clk), .Reset(Reset), .Xc(10'd383), .Yc(10'd67), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[224]) );

cookie ck225 (.Clk(Clk), .Reset(Reset), .Xc(10'd369), .Yc(10'd67), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[225]) );

cookie ck226 (.Clk(Clk), .Reset(Reset), .Xc(10'd355), .Yc(10'd67), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[226]) );

cookie ck227 (.Clk(Clk), .Reset(Reset), .Xc(10'd341), .Yc(10'd67), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[227]) );

cookie ck228 (.Clk(Clk), .Reset(Reset), .Xc(10'd298), .Yc(10'd67), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[228]) );

cookie ck229 (.Clk(Clk), .Reset(Reset), .Xc(10'd283), .Yc(10'd67), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[229]) );

cookie ck230 (.Clk(Clk), .Reset(Reset), .Xc(10'd269), .Yc(10'd67), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[230]) );

cookie ck231 (.Clk(Clk), .Reset(Reset), .Xc(10'd255), .Yc(10'd67), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[231]) );

cookie ck232 (.Clk(Clk), .Reset(Reset), .Xc(10'd241), .Yc(10'd67), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[232]) );

cookie ck233 (.Clk(Clk), .Reset(Reset), .Xc(10'd226), .Yc(10'd67), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[233]) );

cookie ck234 (.Clk(Clk), .Reset(Reset), .Xc(10'd212), .Yc(10'd67), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[234]) );

cookie ck235 (.Clk(Clk), .Reset(Reset), .Xc(10'd198), .Yc(10'd67), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[235]) );

cookie ck236 (.Clk(Clk), .Reset(Reset), .Xc(10'd183), .Yc(10'd67), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[236]) );

cookie ck237 (.Clk(Clk), .Reset(Reset), .Xc(10'd169), .Yc(10'd67), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[237]) );

cookie ck238 (.Clk(Clk), .Reset(Reset), .Xc(10'd155), .Yc(10'd67), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[238]) );

cookie ck239 (.Clk(Clk), .Reset(Reset), .Xc(10'd141), .Yc(10'd67), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[239]) );

cookie ck240 (.Clk(Clk), .Reset(Reset), .Xc(10'd319), .Yc(10'd239), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[240]) );



endmodule

