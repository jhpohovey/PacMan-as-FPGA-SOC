`define COOKIE_COUNT 240

module cookies_wrapper_all (
	input logic Reset,
	input logic Clk,
	input logic [9:0] BallX,
	input logic [9:0] BallY,
	input logic [9:0] Ball_Size,

	output logic [7:0] Total_Score,
	output logic [`COOKIE_COUNT-1:0] Not_ate
);

logic summation_tmp;
reg [`COOKIE_COUNT-1:0] cookie_scores;



integer i;
always_comb begin
	for(i = 0; i < `COOKIE_COUNT; i = i + 1) begin
		summation_tmp += cookie_scores[i];
	end
end


always_ff @ (posedge Clk or posedge Reset)begin
	if (Reset) Total_Score <= 1'b0;
	else Total_Score <= summation_tmp;
end

cookie ck0 (.Clk(Clk), .Reset(Reset), .Xc(10'd498), .Yc(10'd428), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[0]), .Score(cookie_scores[0]) );

cookie ck1 (.Clk(Clk), .Reset(Reset), .Xc(10'd483), .Yc(10'd428), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[1]), .Score(cookie_scores[1]) );

cookie ck2 (.Clk(Clk), .Reset(Reset), .Xc(10'd469), .Yc(10'd428), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[2]), .Score(cookie_scores[2]) );

cookie ck3 (.Clk(Clk), .Reset(Reset), .Xc(10'd455), .Yc(10'd428), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[3]), .Score(cookie_scores[3]) );

cookie ck4 (.Clk(Clk), .Reset(Reset), .Xc(10'd441), .Yc(10'd428), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[4]), .Score(cookie_scores[4]) );

cookie ck5 (.Clk(Clk), .Reset(Reset), .Xc(10'd426), .Yc(10'd428), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[5]), .Score(cookie_scores[5]) );

cookie ck6 (.Clk(Clk), .Reset(Reset), .Xc(10'd412), .Yc(10'd428), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[6]), .Score(cookie_scores[6]) );

cookie ck7 (.Clk(Clk), .Reset(Reset), .Xc(10'd398), .Yc(10'd428), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[7]), .Score(cookie_scores[7]) );

cookie ck8 (.Clk(Clk), .Reset(Reset), .Xc(10'd383), .Yc(10'd428), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[8]), .Score(cookie_scores[8]) );

cookie ck9 (.Clk(Clk), .Reset(Reset), .Xc(10'd369), .Yc(10'd428), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[9]), .Score(cookie_scores[9]) );

cookie ck10 (.Clk(Clk), .Reset(Reset), .Xc(10'd355), .Yc(10'd428), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[10]), .Score(cookie_scores[10]) );

cookie ck11 (.Clk(Clk), .Reset(Reset), .Xc(10'd341), .Yc(10'd428), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[11]), .Score(cookie_scores[11]) );

cookie ck12 (.Clk(Clk), .Reset(Reset), .Xc(10'd326), .Yc(10'd428), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[12]), .Score(cookie_scores[12]) );

cookie ck13 (.Clk(Clk), .Reset(Reset), .Xc(10'd312), .Yc(10'd428), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[13]), .Score(cookie_scores[13]) );

cookie ck14 (.Clk(Clk), .Reset(Reset), .Xc(10'd298), .Yc(10'd428), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[14]), .Score(cookie_scores[14]) );

cookie ck15 (.Clk(Clk), .Reset(Reset), .Xc(10'd283), .Yc(10'd428), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[15]), .Score(cookie_scores[15]) );

cookie ck16 (.Clk(Clk), .Reset(Reset), .Xc(10'd269), .Yc(10'd428), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[16]), .Score(cookie_scores[16]) );

cookie ck17 (.Clk(Clk), .Reset(Reset), .Xc(10'd255), .Yc(10'd428), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[17]), .Score(cookie_scores[17]) );

cookie ck18 (.Clk(Clk), .Reset(Reset), .Xc(10'd241), .Yc(10'd428), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[18]), .Score(cookie_scores[18]) );

cookie ck19 (.Clk(Clk), .Reset(Reset), .Xc(10'd226), .Yc(10'd428), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[19]), .Score(cookie_scores[19]) );

cookie ck20 (.Clk(Clk), .Reset(Reset), .Xc(10'd212), .Yc(10'd428), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[20]), .Score(cookie_scores[20]) );

cookie ck21 (.Clk(Clk), .Reset(Reset), .Xc(10'd198), .Yc(10'd428), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[21]), .Score(cookie_scores[21]) );

cookie ck22 (.Clk(Clk), .Reset(Reset), .Xc(10'd183), .Yc(10'd428), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[22]), .Score(cookie_scores[22]) );

cookie ck23 (.Clk(Clk), .Reset(Reset), .Xc(10'd169), .Yc(10'd428), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[23]), .Score(cookie_scores[23]) );

cookie ck24 (.Clk(Clk), .Reset(Reset), .Xc(10'd155), .Yc(10'd428), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[24]), .Score(cookie_scores[24]) );

cookie ck25 (.Clk(Clk), .Reset(Reset), .Xc(10'd141), .Yc(10'd428), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[25]), .Score(cookie_scores[25]) );

cookie ck26 (.Clk(Clk), .Reset(Reset), .Xc(10'd498), .Yc(10'd415), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[26]), .Score(cookie_scores[26]) );

cookie ck27 (.Clk(Clk), .Reset(Reset), .Xc(10'd341), .Yc(10'd415), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[27]), .Score(cookie_scores[27]) );

cookie ck28 (.Clk(Clk), .Reset(Reset), .Xc(10'd298), .Yc(10'd415), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[28]), .Score(cookie_scores[28]) );

cookie ck29 (.Clk(Clk), .Reset(Reset), .Xc(10'd141), .Yc(10'd415), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[29]), .Score(cookie_scores[29]) );

cookie ck30 (.Clk(Clk), .Reset(Reset), .Xc(10'd498), .Yc(10'd402), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[30]), .Score(cookie_scores[30]) );

cookie ck31 (.Clk(Clk), .Reset(Reset), .Xc(10'd341), .Yc(10'd402), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[31]), .Score(cookie_scores[31]) );

cookie ck32 (.Clk(Clk), .Reset(Reset), .Xc(10'd298), .Yc(10'd402), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[32]), .Score(cookie_scores[32]) );

cookie ck33 (.Clk(Clk), .Reset(Reset), .Xc(10'd141), .Yc(10'd402), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[33]), .Score(cookie_scores[33]) );

cookie ck34 (.Clk(Clk), .Reset(Reset), .Xc(10'd498), .Yc(10'd389), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[34]), .Score(cookie_scores[34]) );

cookie ck35 (.Clk(Clk), .Reset(Reset), .Xc(10'd483), .Yc(10'd389), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[35]), .Score(cookie_scores[35]) );

cookie ck36 (.Clk(Clk), .Reset(Reset), .Xc(10'd469), .Yc(10'd389), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[36]), .Score(cookie_scores[36]) );

cookie ck37 (.Clk(Clk), .Reset(Reset), .Xc(10'd455), .Yc(10'd389), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[37]), .Score(cookie_scores[37]) );

cookie ck38 (.Clk(Clk), .Reset(Reset), .Xc(10'd441), .Yc(10'd389), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[38]), .Score(cookie_scores[38]) );

cookie ck39 (.Clk(Clk), .Reset(Reset), .Xc(10'd426), .Yc(10'd389), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[39]), .Score(cookie_scores[39]) );

cookie ck40 (.Clk(Clk), .Reset(Reset), .Xc(10'd383), .Yc(10'd389), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[40]), .Score(cookie_scores[40]) );

cookie ck41 (.Clk(Clk), .Reset(Reset), .Xc(10'd369), .Yc(10'd389), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[41]), .Score(cookie_scores[41]) );

cookie ck42 (.Clk(Clk), .Reset(Reset), .Xc(10'd355), .Yc(10'd389), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[42]), .Score(cookie_scores[42]) );

cookie ck43 (.Clk(Clk), .Reset(Reset), .Xc(10'd341), .Yc(10'd389), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[43]), .Score(cookie_scores[43]) );

cookie ck44 (.Clk(Clk), .Reset(Reset), .Xc(10'd298), .Yc(10'd389), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[44]), .Score(cookie_scores[44]) );

cookie ck45 (.Clk(Clk), .Reset(Reset), .Xc(10'd283), .Yc(10'd389), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[45]), .Score(cookie_scores[45]) );

cookie ck46 (.Clk(Clk), .Reset(Reset), .Xc(10'd269), .Yc(10'd389), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[46]), .Score(cookie_scores[46]) );

cookie ck47 (.Clk(Clk), .Reset(Reset), .Xc(10'd255), .Yc(10'd389), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[47]), .Score(cookie_scores[47]) );

cookie ck48 (.Clk(Clk), .Reset(Reset), .Xc(10'd212), .Yc(10'd389), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[48]), .Score(cookie_scores[48]) );

cookie ck49 (.Clk(Clk), .Reset(Reset), .Xc(10'd198), .Yc(10'd389), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[49]), .Score(cookie_scores[49]) );

cookie ck50 (.Clk(Clk), .Reset(Reset), .Xc(10'd183), .Yc(10'd389), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[50]), .Score(cookie_scores[50]) );

cookie ck51 (.Clk(Clk), .Reset(Reset), .Xc(10'd169), .Yc(10'd389), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[51]), .Score(cookie_scores[51]) );

cookie ck52 (.Clk(Clk), .Reset(Reset), .Xc(10'd155), .Yc(10'd389), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[52]), .Score(cookie_scores[52]) );

cookie ck53 (.Clk(Clk), .Reset(Reset), .Xc(10'd141), .Yc(10'd389), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[53]), .Score(cookie_scores[53]) );

cookie ck54 (.Clk(Clk), .Reset(Reset), .Xc(10'd469), .Yc(10'd376), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[54]), .Score(cookie_scores[54]) );

cookie ck55 (.Clk(Clk), .Reset(Reset), .Xc(10'd426), .Yc(10'd376), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[55]), .Score(cookie_scores[55]) );

cookie ck56 (.Clk(Clk), .Reset(Reset), .Xc(10'd383), .Yc(10'd376), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[56]), .Score(cookie_scores[56]) );

cookie ck57 (.Clk(Clk), .Reset(Reset), .Xc(10'd255), .Yc(10'd376), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[57]), .Score(cookie_scores[57]) );

cookie ck58 (.Clk(Clk), .Reset(Reset), .Xc(10'd212), .Yc(10'd376), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[58]), .Score(cookie_scores[58]) );

cookie ck59 (.Clk(Clk), .Reset(Reset), .Xc(10'd169), .Yc(10'd376), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[59]), .Score(cookie_scores[59]) );

cookie ck60 (.Clk(Clk), .Reset(Reset), .Xc(10'd469), .Yc(10'd364), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[60]), .Score(cookie_scores[60]) );

cookie ck61 (.Clk(Clk), .Reset(Reset), .Xc(10'd426), .Yc(10'd364), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[61]), .Score(cookie_scores[61]) );

cookie ck62 (.Clk(Clk), .Reset(Reset), .Xc(10'd383), .Yc(10'd364), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[62]), .Score(cookie_scores[62]) );

cookie ck63 (.Clk(Clk), .Reset(Reset), .Xc(10'd255), .Yc(10'd364), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[63]), .Score(cookie_scores[63]) );

cookie ck64 (.Clk(Clk), .Reset(Reset), .Xc(10'd212), .Yc(10'd364), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[64]), .Score(cookie_scores[64]) );

cookie ck65 (.Clk(Clk), .Reset(Reset), .Xc(10'd169), .Yc(10'd364), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[65]), .Score(cookie_scores[65]) );

cookie ck66 (.Clk(Clk), .Reset(Reset), .Xc(10'd483), .Yc(10'd351), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[66]), .Score(cookie_scores[66]) );

cookie ck67 (.Clk(Clk), .Reset(Reset), .Xc(10'd469), .Yc(10'd351), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[67]), .Score(cookie_scores[67]) );

cookie ck68 (.Clk(Clk), .Reset(Reset), .Xc(10'd426), .Yc(10'd351), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[68]), .Score(cookie_scores[68]) );

cookie ck69 (.Clk(Clk), .Reset(Reset), .Xc(10'd412), .Yc(10'd351), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[69]), .Score(cookie_scores[69]) );

cookie ck70 (.Clk(Clk), .Reset(Reset), .Xc(10'd398), .Yc(10'd351), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[70]), .Score(cookie_scores[70]) );

cookie ck71 (.Clk(Clk), .Reset(Reset), .Xc(10'd383), .Yc(10'd351), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[71]), .Score(cookie_scores[71]) );

cookie ck72 (.Clk(Clk), .Reset(Reset), .Xc(10'd369), .Yc(10'd351), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[72]), .Score(cookie_scores[72]) );

cookie ck73 (.Clk(Clk), .Reset(Reset), .Xc(10'd355), .Yc(10'd351), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[73]), .Score(cookie_scores[73]) );

cookie ck74 (.Clk(Clk), .Reset(Reset), .Xc(10'd341), .Yc(10'd351), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[74]), .Score(cookie_scores[74]) );

cookie ck75 (.Clk(Clk), .Reset(Reset), .Xc(10'd298), .Yc(10'd351), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[75]), .Score(cookie_scores[75]) );

cookie ck76 (.Clk(Clk), .Reset(Reset), .Xc(10'd283), .Yc(10'd351), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[76]), .Score(cookie_scores[76]) );

cookie ck77 (.Clk(Clk), .Reset(Reset), .Xc(10'd269), .Yc(10'd351), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[77]), .Score(cookie_scores[77]) );

cookie ck78 (.Clk(Clk), .Reset(Reset), .Xc(10'd255), .Yc(10'd351), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[78]), .Score(cookie_scores[78]) );

cookie ck79 (.Clk(Clk), .Reset(Reset), .Xc(10'd241), .Yc(10'd351), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[79]), .Score(cookie_scores[79]) );

cookie ck80 (.Clk(Clk), .Reset(Reset), .Xc(10'd226), .Yc(10'd351), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[80]), .Score(cookie_scores[80]) );

cookie ck81 (.Clk(Clk), .Reset(Reset), .Xc(10'd212), .Yc(10'd351), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[81]), .Score(cookie_scores[81]) );

cookie ck82 (.Clk(Clk), .Reset(Reset), .Xc(10'd169), .Yc(10'd351), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[82]), .Score(cookie_scores[82]) );

cookie ck83 (.Clk(Clk), .Reset(Reset), .Xc(10'd155), .Yc(10'd351), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[83]), .Score(cookie_scores[83]) );

cookie ck84 (.Clk(Clk), .Reset(Reset), .Xc(10'd498), .Yc(10'd338), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[84]), .Score(cookie_scores[84]) );

cookie ck85 (.Clk(Clk), .Reset(Reset), .Xc(10'd426), .Yc(10'd338), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[85]), .Score(cookie_scores[85]) );

cookie ck86 (.Clk(Clk), .Reset(Reset), .Xc(10'd341), .Yc(10'd338), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[86]), .Score(cookie_scores[86]) );

cookie ck87 (.Clk(Clk), .Reset(Reset), .Xc(10'd298), .Yc(10'd338), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[87]), .Score(cookie_scores[87]) );

cookie ck88 (.Clk(Clk), .Reset(Reset), .Xc(10'd212), .Yc(10'd338), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[88]), .Score(cookie_scores[88]) );

cookie ck89 (.Clk(Clk), .Reset(Reset), .Xc(10'd141), .Yc(10'd338), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[89]), .Score(cookie_scores[89]) );

cookie ck90 (.Clk(Clk), .Reset(Reset), .Xc(10'd498), .Yc(10'd325), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[90]), .Score(cookie_scores[90]) );

cookie ck91 (.Clk(Clk), .Reset(Reset), .Xc(10'd426), .Yc(10'd325), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[91]), .Score(cookie_scores[91]) );

cookie ck92 (.Clk(Clk), .Reset(Reset), .Xc(10'd341), .Yc(10'd325), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[92]), .Score(cookie_scores[92]) );

cookie ck93 (.Clk(Clk), .Reset(Reset), .Xc(10'd298), .Yc(10'd325), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[93]), .Score(cookie_scores[93]) );

cookie ck94 (.Clk(Clk), .Reset(Reset), .Xc(10'd212), .Yc(10'd325), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[94]), .Score(cookie_scores[94]) );

cookie ck95 (.Clk(Clk), .Reset(Reset), .Xc(10'd141), .Yc(10'd325), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[95]), .Score(cookie_scores[95]) );

cookie ck96 (.Clk(Clk), .Reset(Reset), .Xc(10'd498), .Yc(10'd312), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[96]), .Score(cookie_scores[96]) );

cookie ck97 (.Clk(Clk), .Reset(Reset), .Xc(10'd483), .Yc(10'd312), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[97]), .Score(cookie_scores[97]) );

cookie ck98 (.Clk(Clk), .Reset(Reset), .Xc(10'd469), .Yc(10'd312), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[98]), .Score(cookie_scores[98]) );

cookie ck99 (.Clk(Clk), .Reset(Reset), .Xc(10'd455), .Yc(10'd312), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[99]), .Score(cookie_scores[99]) );

cookie ck100 (.Clk(Clk), .Reset(Reset), .Xc(10'd441), .Yc(10'd312), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[100]), .Score(cookie_scores[100]) );

cookie ck101 (.Clk(Clk), .Reset(Reset), .Xc(10'd426), .Yc(10'd312), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[101]), .Score(cookie_scores[101]) );

cookie ck102 (.Clk(Clk), .Reset(Reset), .Xc(10'd412), .Yc(10'd312), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[102]), .Score(cookie_scores[102]) );

cookie ck103 (.Clk(Clk), .Reset(Reset), .Xc(10'd398), .Yc(10'd312), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[103]), .Score(cookie_scores[103]) );

cookie ck104 (.Clk(Clk), .Reset(Reset), .Xc(10'd383), .Yc(10'd312), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[104]), .Score(cookie_scores[104]) );

cookie ck105 (.Clk(Clk), .Reset(Reset), .Xc(10'd369), .Yc(10'd312), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[105]), .Score(cookie_scores[105]) );

cookie ck106 (.Clk(Clk), .Reset(Reset), .Xc(10'd355), .Yc(10'd312), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[106]), .Score(cookie_scores[106]) );

cookie ck107 (.Clk(Clk), .Reset(Reset), .Xc(10'd341), .Yc(10'd312), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[107]), .Score(cookie_scores[107]) );

cookie ck108 (.Clk(Clk), .Reset(Reset), .Xc(10'd298), .Yc(10'd312), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[108]), .Score(cookie_scores[108]) );

cookie ck109 (.Clk(Clk), .Reset(Reset), .Xc(10'd283), .Yc(10'd312), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[109]), .Score(cookie_scores[109]) );

cookie ck110 (.Clk(Clk), .Reset(Reset), .Xc(10'd269), .Yc(10'd312), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[110]), .Score(cookie_scores[110]) );

cookie ck111 (.Clk(Clk), .Reset(Reset), .Xc(10'd255), .Yc(10'd312), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[111]), .Score(cookie_scores[111]) );

cookie ck112 (.Clk(Clk), .Reset(Reset), .Xc(10'd241), .Yc(10'd312), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[112]), .Score(cookie_scores[112]) );

cookie ck113 (.Clk(Clk), .Reset(Reset), .Xc(10'd226), .Yc(10'd312), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[113]), .Score(cookie_scores[113]) );

cookie ck114 (.Clk(Clk), .Reset(Reset), .Xc(10'd212), .Yc(10'd312), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[114]), .Score(cookie_scores[114]) );

cookie ck115 (.Clk(Clk), .Reset(Reset), .Xc(10'd198), .Yc(10'd312), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[115]), .Score(cookie_scores[115]) );

cookie ck116 (.Clk(Clk), .Reset(Reset), .Xc(10'd183), .Yc(10'd312), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[116]), .Score(cookie_scores[116]) );

cookie ck117 (.Clk(Clk), .Reset(Reset), .Xc(10'd169), .Yc(10'd312), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[117]), .Score(cookie_scores[117]) );

cookie ck118 (.Clk(Clk), .Reset(Reset), .Xc(10'd155), .Yc(10'd312), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[118]), .Score(cookie_scores[118]) );

cookie ck119 (.Clk(Clk), .Reset(Reset), .Xc(10'd141), .Yc(10'd312), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[119]), .Score(cookie_scores[119]) );

cookie ck120 (.Clk(Clk), .Reset(Reset), .Xc(10'd426), .Yc(10'd299), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[120]), .Score(cookie_scores[120]) );

cookie ck121 (.Clk(Clk), .Reset(Reset), .Xc(10'd212), .Yc(10'd299), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[121]), .Score(cookie_scores[121]) );

cookie ck122 (.Clk(Clk), .Reset(Reset), .Xc(10'd426), .Yc(10'd286), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[122]), .Score(cookie_scores[122]) );

cookie ck123 (.Clk(Clk), .Reset(Reset), .Xc(10'd212), .Yc(10'd286), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[123]), .Score(cookie_scores[123]) );

cookie ck124 (.Clk(Clk), .Reset(Reset), .Xc(10'd426), .Yc(10'd273), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[124]), .Score(cookie_scores[124]) );

cookie ck125 (.Clk(Clk), .Reset(Reset), .Xc(10'd212), .Yc(10'd273), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[125]), .Score(cookie_scores[125]) );

cookie ck126 (.Clk(Clk), .Reset(Reset), .Xc(10'd426), .Yc(10'd260), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[126]), .Score(cookie_scores[126]) );

cookie ck127 (.Clk(Clk), .Reset(Reset), .Xc(10'd212), .Yc(10'd260), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[127]), .Score(cookie_scores[127]) );

cookie ck128 (.Clk(Clk), .Reset(Reset), .Xc(10'd426), .Yc(10'd247), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[128]), .Score(cookie_scores[128]) );

cookie ck129 (.Clk(Clk), .Reset(Reset), .Xc(10'd212), .Yc(10'd247), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[129]), .Score(cookie_scores[129]) );

cookie ck130 (.Clk(Clk), .Reset(Reset), .Xc(10'd426), .Yc(10'd234), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[130]), .Score(cookie_scores[130]) );

cookie ck131 (.Clk(Clk), .Reset(Reset), .Xc(10'd212), .Yc(10'd234), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[131]), .Score(cookie_scores[131]) );

cookie ck132 (.Clk(Clk), .Reset(Reset), .Xc(10'd426), .Yc(10'd222), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[132]), .Score(cookie_scores[132]) );

cookie ck133 (.Clk(Clk), .Reset(Reset), .Xc(10'd212), .Yc(10'd222), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[133]), .Score(cookie_scores[133]) );

cookie ck134 (.Clk(Clk), .Reset(Reset), .Xc(10'd426), .Yc(10'd209), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[134]), .Score(cookie_scores[134]) );

cookie ck135 (.Clk(Clk), .Reset(Reset), .Xc(10'd212), .Yc(10'd209), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[135]), .Score(cookie_scores[135]) );

cookie ck136 (.Clk(Clk), .Reset(Reset), .Xc(10'd426), .Yc(10'd196), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[136]), .Score(cookie_scores[136]) );

cookie ck137 (.Clk(Clk), .Reset(Reset), .Xc(10'd212), .Yc(10'd196), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[137]), .Score(cookie_scores[137]) );

cookie ck138 (.Clk(Clk), .Reset(Reset), .Xc(10'd426), .Yc(10'd183), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[138]), .Score(cookie_scores[138]) );

cookie ck139 (.Clk(Clk), .Reset(Reset), .Xc(10'd212), .Yc(10'd183), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[139]), .Score(cookie_scores[139]) );

cookie ck140 (.Clk(Clk), .Reset(Reset), .Xc(10'd426), .Yc(10'd170), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[140]), .Score(cookie_scores[140]) );

cookie ck141 (.Clk(Clk), .Reset(Reset), .Xc(10'd212), .Yc(10'd170), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[141]), .Score(cookie_scores[141]) );

cookie ck142 (.Clk(Clk), .Reset(Reset), .Xc(10'd498), .Yc(10'd157), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[142]), .Score(cookie_scores[142]) );

cookie ck143 (.Clk(Clk), .Reset(Reset), .Xc(10'd483), .Yc(10'd157), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[143]), .Score(cookie_scores[143]) );

cookie ck144 (.Clk(Clk), .Reset(Reset), .Xc(10'd469), .Yc(10'd157), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[144]), .Score(cookie_scores[144]) );

cookie ck145 (.Clk(Clk), .Reset(Reset), .Xc(10'd455), .Yc(10'd157), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[145]), .Score(cookie_scores[145]) );

cookie ck146 (.Clk(Clk), .Reset(Reset), .Xc(10'd441), .Yc(10'd157), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[146]), .Score(cookie_scores[146]) );

cookie ck147 (.Clk(Clk), .Reset(Reset), .Xc(10'd426), .Yc(10'd157), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[147]), .Score(cookie_scores[147]) );

cookie ck148 (.Clk(Clk), .Reset(Reset), .Xc(10'd383), .Yc(10'd157), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[148]), .Score(cookie_scores[148]) );

cookie ck149 (.Clk(Clk), .Reset(Reset), .Xc(10'd369), .Yc(10'd157), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[149]), .Score(cookie_scores[149]) );

cookie ck150 (.Clk(Clk), .Reset(Reset), .Xc(10'd355), .Yc(10'd157), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[150]), .Score(cookie_scores[150]) );

cookie ck151 (.Clk(Clk), .Reset(Reset), .Xc(10'd341), .Yc(10'd157), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[151]), .Score(cookie_scores[151]) );

cookie ck152 (.Clk(Clk), .Reset(Reset), .Xc(10'd298), .Yc(10'd157), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[152]), .Score(cookie_scores[152]) );

cookie ck153 (.Clk(Clk), .Reset(Reset), .Xc(10'd283), .Yc(10'd157), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[153]), .Score(cookie_scores[153]) );

cookie ck154 (.Clk(Clk), .Reset(Reset), .Xc(10'd269), .Yc(10'd157), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[154]), .Score(cookie_scores[154]) );

cookie ck155 (.Clk(Clk), .Reset(Reset), .Xc(10'd255), .Yc(10'd157), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[155]), .Score(cookie_scores[155]) );

cookie ck156 (.Clk(Clk), .Reset(Reset), .Xc(10'd212), .Yc(10'd157), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[156]), .Score(cookie_scores[156]) );

cookie ck157 (.Clk(Clk), .Reset(Reset), .Xc(10'd198), .Yc(10'd157), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[157]), .Score(cookie_scores[157]) );

cookie ck158 (.Clk(Clk), .Reset(Reset), .Xc(10'd183), .Yc(10'd157), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[158]), .Score(cookie_scores[158]) );

cookie ck159 (.Clk(Clk), .Reset(Reset), .Xc(10'd169), .Yc(10'd157), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[159]), .Score(cookie_scores[159]) );

cookie ck160 (.Clk(Clk), .Reset(Reset), .Xc(10'd155), .Yc(10'd157), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[160]), .Score(cookie_scores[160]) );

cookie ck161 (.Clk(Clk), .Reset(Reset), .Xc(10'd141), .Yc(10'd157), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[161]), .Score(cookie_scores[161]) );

cookie ck162 (.Clk(Clk), .Reset(Reset), .Xc(10'd498), .Yc(10'd144), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[162]), .Score(cookie_scores[162]) );

cookie ck163 (.Clk(Clk), .Reset(Reset), .Xc(10'd426), .Yc(10'd144), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[163]), .Score(cookie_scores[163]) );

cookie ck164 (.Clk(Clk), .Reset(Reset), .Xc(10'd383), .Yc(10'd144), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[164]), .Score(cookie_scores[164]) );

cookie ck165 (.Clk(Clk), .Reset(Reset), .Xc(10'd255), .Yc(10'd144), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[165]), .Score(cookie_scores[165]) );

cookie ck166 (.Clk(Clk), .Reset(Reset), .Xc(10'd212), .Yc(10'd144), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[166]), .Score(cookie_scores[166]) );

cookie ck167 (.Clk(Clk), .Reset(Reset), .Xc(10'd141), .Yc(10'd144), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[167]), .Score(cookie_scores[167]) );

cookie ck168 (.Clk(Clk), .Reset(Reset), .Xc(10'd498), .Yc(10'd131), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[168]), .Score(cookie_scores[168]) );

cookie ck169 (.Clk(Clk), .Reset(Reset), .Xc(10'd426), .Yc(10'd131), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[169]), .Score(cookie_scores[169]) );

cookie ck170 (.Clk(Clk), .Reset(Reset), .Xc(10'd383), .Yc(10'd131), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[170]), .Score(cookie_scores[170]) );

cookie ck171 (.Clk(Clk), .Reset(Reset), .Xc(10'd255), .Yc(10'd131), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[171]), .Score(cookie_scores[171]) );

cookie ck172 (.Clk(Clk), .Reset(Reset), .Xc(10'd212), .Yc(10'd131), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[172]), .Score(cookie_scores[172]) );

cookie ck173 (.Clk(Clk), .Reset(Reset), .Xc(10'd141), .Yc(10'd131), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[173]), .Score(cookie_scores[173]) );

cookie ck174 (.Clk(Clk), .Reset(Reset), .Xc(10'd498), .Yc(10'd118), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[174]), .Score(cookie_scores[174]) );

cookie ck175 (.Clk(Clk), .Reset(Reset), .Xc(10'd483), .Yc(10'd118), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[175]), .Score(cookie_scores[175]) );

cookie ck176 (.Clk(Clk), .Reset(Reset), .Xc(10'd469), .Yc(10'd118), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[176]), .Score(cookie_scores[176]) );

cookie ck177 (.Clk(Clk), .Reset(Reset), .Xc(10'd455), .Yc(10'd118), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[177]), .Score(cookie_scores[177]) );

cookie ck178 (.Clk(Clk), .Reset(Reset), .Xc(10'd441), .Yc(10'd118), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[178]), .Score(cookie_scores[178]) );

cookie ck179 (.Clk(Clk), .Reset(Reset), .Xc(10'd426), .Yc(10'd118), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[179]), .Score(cookie_scores[179]) );

cookie ck180 (.Clk(Clk), .Reset(Reset), .Xc(10'd412), .Yc(10'd118), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[180]), .Score(cookie_scores[180]) );

cookie ck181 (.Clk(Clk), .Reset(Reset), .Xc(10'd398), .Yc(10'd118), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[181]), .Score(cookie_scores[181]) );

cookie ck182 (.Clk(Clk), .Reset(Reset), .Xc(10'd383), .Yc(10'd118), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[182]), .Score(cookie_scores[182]) );

cookie ck183 (.Clk(Clk), .Reset(Reset), .Xc(10'd369), .Yc(10'd118), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[183]), .Score(cookie_scores[183]) );

cookie ck184 (.Clk(Clk), .Reset(Reset), .Xc(10'd355), .Yc(10'd118), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[184]), .Score(cookie_scores[184]) );

cookie ck185 (.Clk(Clk), .Reset(Reset), .Xc(10'd341), .Yc(10'd118), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[185]), .Score(cookie_scores[185]) );

cookie ck186 (.Clk(Clk), .Reset(Reset), .Xc(10'd326), .Yc(10'd118), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[186]), .Score(cookie_scores[186]) );

cookie ck187 (.Clk(Clk), .Reset(Reset), .Xc(10'd312), .Yc(10'd118), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[187]), .Score(cookie_scores[187]) );

cookie ck188 (.Clk(Clk), .Reset(Reset), .Xc(10'd298), .Yc(10'd118), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[188]), .Score(cookie_scores[188]) );

cookie ck189 (.Clk(Clk), .Reset(Reset), .Xc(10'd283), .Yc(10'd118), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[189]), .Score(cookie_scores[189]) );

cookie ck190 (.Clk(Clk), .Reset(Reset), .Xc(10'd269), .Yc(10'd118), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[190]), .Score(cookie_scores[190]) );

cookie ck191 (.Clk(Clk), .Reset(Reset), .Xc(10'd255), .Yc(10'd118), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[191]), .Score(cookie_scores[191]) );

cookie ck192 (.Clk(Clk), .Reset(Reset), .Xc(10'd241), .Yc(10'd118), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[192]), .Score(cookie_scores[192]) );

cookie ck193 (.Clk(Clk), .Reset(Reset), .Xc(10'd226), .Yc(10'd118), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[193]), .Score(cookie_scores[193]) );

cookie ck194 (.Clk(Clk), .Reset(Reset), .Xc(10'd212), .Yc(10'd118), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[194]), .Score(cookie_scores[194]) );

cookie ck195 (.Clk(Clk), .Reset(Reset), .Xc(10'd198), .Yc(10'd118), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[195]), .Score(cookie_scores[195]) );

cookie ck196 (.Clk(Clk), .Reset(Reset), .Xc(10'd183), .Yc(10'd118), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[196]), .Score(cookie_scores[196]) );

cookie ck197 (.Clk(Clk), .Reset(Reset), .Xc(10'd169), .Yc(10'd118), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[197]), .Score(cookie_scores[197]) );

cookie ck198 (.Clk(Clk), .Reset(Reset), .Xc(10'd155), .Yc(10'd118), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[198]), .Score(cookie_scores[198]) );

cookie ck199 (.Clk(Clk), .Reset(Reset), .Xc(10'd141), .Yc(10'd118), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[199]), .Score(cookie_scores[199]) );

cookie ck200 (.Clk(Clk), .Reset(Reset), .Xc(10'd498), .Yc(10'd105), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[200]), .Score(cookie_scores[200]) );

cookie ck201 (.Clk(Clk), .Reset(Reset), .Xc(10'd341), .Yc(10'd105), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[201]), .Score(cookie_scores[201]) );

cookie ck202 (.Clk(Clk), .Reset(Reset), .Xc(10'd298), .Yc(10'd105), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[202]), .Score(cookie_scores[202]) );

cookie ck203 (.Clk(Clk), .Reset(Reset), .Xc(10'd141), .Yc(10'd105), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[203]), .Score(cookie_scores[203]) );

cookie ck204 (.Clk(Clk), .Reset(Reset), .Xc(10'd426), .Yc(10'd105), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[204]), .Score(cookie_scores[204]) );

cookie ck205 (.Clk(Clk), .Reset(Reset), .Xc(10'd212), .Yc(10'd105), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[205]), .Score(cookie_scores[205]) );

cookie ck206 (.Clk(Clk), .Reset(Reset), .Xc(10'd426), .Yc(10'd93), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[206]), .Score(cookie_scores[206]) );

cookie ck207 (.Clk(Clk), .Reset(Reset), .Xc(10'd341), .Yc(10'd93), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[207]), .Score(cookie_scores[207]) );

cookie ck208 (.Clk(Clk), .Reset(Reset), .Xc(10'd298), .Yc(10'd93), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[208]), .Score(cookie_scores[208]) );

cookie ck209 (.Clk(Clk), .Reset(Reset), .Xc(10'd212), .Yc(10'd93), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[209]), .Score(cookie_scores[209]) );

cookie ck210 (.Clk(Clk), .Reset(Reset), .Xc(10'd498), .Yc(10'd80), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[210]), .Score(cookie_scores[210]) );

cookie ck211 (.Clk(Clk), .Reset(Reset), .Xc(10'd426), .Yc(10'd80), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[211]), .Score(cookie_scores[211]) );

cookie ck212 (.Clk(Clk), .Reset(Reset), .Xc(10'd341), .Yc(10'd80), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[212]), .Score(cookie_scores[212]) );

cookie ck213 (.Clk(Clk), .Reset(Reset), .Xc(10'd298), .Yc(10'd80), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[213]), .Score(cookie_scores[213]) );

cookie ck214 (.Clk(Clk), .Reset(Reset), .Xc(10'd212), .Yc(10'd80), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[214]), .Score(cookie_scores[214]) );

cookie ck215 (.Clk(Clk), .Reset(Reset), .Xc(10'd141), .Yc(10'd80), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[215]), .Score(cookie_scores[215]) );

cookie ck216 (.Clk(Clk), .Reset(Reset), .Xc(10'd498), .Yc(10'd67), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[216]), .Score(cookie_scores[216]) );

cookie ck217 (.Clk(Clk), .Reset(Reset), .Xc(10'd483), .Yc(10'd67), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[217]), .Score(cookie_scores[217]) );

cookie ck218 (.Clk(Clk), .Reset(Reset), .Xc(10'd469), .Yc(10'd67), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[218]), .Score(cookie_scores[218]) );

cookie ck219 (.Clk(Clk), .Reset(Reset), .Xc(10'd455), .Yc(10'd67), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[219]), .Score(cookie_scores[219]) );

cookie ck220 (.Clk(Clk), .Reset(Reset), .Xc(10'd441), .Yc(10'd67), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[220]), .Score(cookie_scores[220]) );

cookie ck221 (.Clk(Clk), .Reset(Reset), .Xc(10'd426), .Yc(10'd67), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[221]), .Score(cookie_scores[221]) );

cookie ck222 (.Clk(Clk), .Reset(Reset), .Xc(10'd412), .Yc(10'd67), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[222]), .Score(cookie_scores[222]) );

cookie ck223 (.Clk(Clk), .Reset(Reset), .Xc(10'd398), .Yc(10'd67), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[223]), .Score(cookie_scores[223]) );

cookie ck224 (.Clk(Clk), .Reset(Reset), .Xc(10'd383), .Yc(10'd67), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[224]), .Score(cookie_scores[224]) );

cookie ck225 (.Clk(Clk), .Reset(Reset), .Xc(10'd369), .Yc(10'd67), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[225]), .Score(cookie_scores[225]) );

cookie ck226 (.Clk(Clk), .Reset(Reset), .Xc(10'd355), .Yc(10'd67), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[226]), .Score(cookie_scores[226]) );

cookie ck227 (.Clk(Clk), .Reset(Reset), .Xc(10'd341), .Yc(10'd67), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[227]), .Score(cookie_scores[227]) );

cookie ck228 (.Clk(Clk), .Reset(Reset), .Xc(10'd298), .Yc(10'd67), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[228]), .Score(cookie_scores[228]) );

cookie ck229 (.Clk(Clk), .Reset(Reset), .Xc(10'd283), .Yc(10'd67), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[229]), .Score(cookie_scores[229]) );

cookie ck230 (.Clk(Clk), .Reset(Reset), .Xc(10'd269), .Yc(10'd67), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[230]), .Score(cookie_scores[230]) );

cookie ck231 (.Clk(Clk), .Reset(Reset), .Xc(10'd255), .Yc(10'd67), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[231]), .Score(cookie_scores[231]) );

cookie ck232 (.Clk(Clk), .Reset(Reset), .Xc(10'd241), .Yc(10'd67), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[232]), .Score(cookie_scores[232]) );

cookie ck233 (.Clk(Clk), .Reset(Reset), .Xc(10'd226), .Yc(10'd67), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[233]), .Score(cookie_scores[233]) );

cookie ck234 (.Clk(Clk), .Reset(Reset), .Xc(10'd212), .Yc(10'd67), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[234]), .Score(cookie_scores[234]) );

cookie ck235 (.Clk(Clk), .Reset(Reset), .Xc(10'd198), .Yc(10'd67), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[235]), .Score(cookie_scores[235]) );

cookie ck236 (.Clk(Clk), .Reset(Reset), .Xc(10'd183), .Yc(10'd67), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[236]), .Score(cookie_scores[236]) );

cookie ck237 (.Clk(Clk), .Reset(Reset), .Xc(10'd169), .Yc(10'd67), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[237]), .Score(cookie_scores[237]) );

cookie ck238 (.Clk(Clk), .Reset(Reset), .Xc(10'd155), .Yc(10'd67), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[238]), .Score(cookie_scores[238]) );

cookie ck239 (.Clk(Clk), .Reset(Reset), .Xc(10'd141), .Yc(10'd67), .Xp(BallX), .Yp(BallY), .Sizep(Ball_Size), .Not_ate(Not_ate[239]), .Score(cookie_scores[239]) );



endmodule

