//module game_end_rom (
//	input [18:0] read_address,
//	input Clk,
//
////	output logic [639:0] data_Out
//	output logic [3:0] data_Out
//
//);
//
//	// mem has width of 128 bits and a total of 256 addresses
////	logic [287:0] mem [0:255];
//	logic [3:0] mem [32768];
//	
//	initial
//	begin
//		 $readmemh("gameover.txt", mem);
//	end
//
//
//	always_ff @ (posedge Clk) begin
//		data_Out<= mem[read_address];
//	end
//
//endmodule
