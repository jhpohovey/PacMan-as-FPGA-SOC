if (DrawY == Y_Pos && DrawX == X_Pos) pixel <=12'h4ff;
if (DrawY == Y_Pos + 0 && DrawX == X_Pos + 1) pixel <=12'h4ff;
if (DrawY == Y_Pos + 0 && DrawX == X_Pos + 2) pixel <=12'h4ff;
if (DrawY == Y_Pos + 0 && DrawX == X_Pos + 3) pixel <=12'h4ff;
if (DrawY == Y_Pos + 0 && DrawX == X_Pos + 4) pixel <=12'h4ff;
if (DrawY == Y_Pos + 0 && DrawX == X_Pos + 5) pixel <=12'h4ff;
if (DrawY == Y_Pos + 0 && DrawX == X_Pos + 6) pixel <= 12'h73f;
if (DrawY == Y_Pos + 0 && DrawX == X_Pos + 7) pixel <=12'h4ff;
if (DrawY == Y_Pos + 0 && DrawX == X_Pos + 8) pixel <=12'h4ff;
if (DrawY == Y_Pos + 0 && DrawX == X_Pos + 9) pixel <=12'h4ff;
if (DrawY == Y_Pos + 0 && DrawX == X_Pos + 10) pixel <= 12'h73f;
if (DrawY == Y_Pos + 0 && DrawX == X_Pos + 11) pixel <= 12'h73f;
if (DrawY == Y_Pos + 0 && DrawX == X_Pos + 12) pixel <=12'h4ff;
if (DrawY == Y_Pos + 0 && DrawX == X_Pos + 13) pixel <=12'h4ff;
if (DrawY == Y_Pos + 0 && DrawX == X_Pos + 14) pixel <=12'h4ff;
if (DrawY == Y_Pos + 0 && DrawX == X_Pos + 15) pixel <=12'h4ff;
if (DrawY == Y_Pos + 1 && DrawX == X_Pos + 0) pixel <=12'h4ff;
if (DrawY == Y_Pos + 1 && DrawX == X_Pos + 1) pixel <=12'h4ff;
if (DrawY == Y_Pos + 1 && DrawX == X_Pos + 2) pixel <=12'h4ff;
if (DrawY == Y_Pos + 1 && DrawX == X_Pos + 3) pixel <=12'h4ff;
if (DrawY == Y_Pos + 1 && DrawX == X_Pos + 4) pixel <= 12'h73f;
if (DrawY == Y_Pos + 1 && DrawX == X_Pos + 5) pixel <= 12'h73f;
if (DrawY == Y_Pos + 1 && DrawX == X_Pos + 6) pixel <=12'h4ff;
if (DrawY == Y_Pos + 1 && DrawX == X_Pos + 7) pixel <= 12'h73f;
if (DrawY == Y_Pos + 1 && DrawX == X_Pos + 8) pixel <= 12'h73f;
if (DrawY == Y_Pos + 1 && DrawX == X_Pos + 9) pixel <= 12'h97d;
if (DrawY == Y_Pos + 1 && DrawX == X_Pos + 10) pixel <= 12'h73f;
if (DrawY == Y_Pos + 1 && DrawX == X_Pos + 11) pixel <=12'h4ff;
if (DrawY == Y_Pos + 1 && DrawX == X_Pos + 12) pixel <= 12'h73f;
if (DrawY == Y_Pos + 1 && DrawX == X_Pos + 13) pixel <=12'h4ff;
if (DrawY == Y_Pos + 1 && DrawX == X_Pos + 14) pixel <= 12'h73f;
if (DrawY == Y_Pos + 1 && DrawX == X_Pos + 15) pixel <=12'h4ff;
if (DrawY == Y_Pos + 2 && DrawX == X_Pos + 0) pixel <= 12'h73f;
if (DrawY == Y_Pos + 2 && DrawX == X_Pos + 1) pixel <=12'h4ff;
if (DrawY == Y_Pos + 2 && DrawX == X_Pos + 2) pixel <=12'h4ff;
if (DrawY == Y_Pos + 2 && DrawX == X_Pos + 3) pixel <= 12'h73f;
if (DrawY == Y_Pos + 2 && DrawX == X_Pos + 4) pixel <=12'h4ff;
if (DrawY == Y_Pos + 2 && DrawX == X_Pos + 5) pixel <= 12'h73f;
if (DrawY == Y_Pos + 2 && DrawX == X_Pos + 6) pixel <= 12'h97d;
if (DrawY == Y_Pos + 2 && DrawX == X_Pos + 7) pixel <= 12'h73f;
if (DrawY == Y_Pos + 2 && DrawX == X_Pos + 8) pixel <=12'h4ff;
if (DrawY == Y_Pos + 2 && DrawX == X_Pos + 9) pixel <= 12'h97d;
if (DrawY == Y_Pos + 2 && DrawX == X_Pos + 10) pixel <=12'h4ff;
if (DrawY == Y_Pos + 2 && DrawX == X_Pos + 11) pixel <= 12'h73f;
if (DrawY == Y_Pos + 2 && DrawX == X_Pos + 12) pixel <= 12'h73f;
if (DrawY == Y_Pos + 2 && DrawX == X_Pos + 13) pixel <=12'h4ff;
if (DrawY == Y_Pos + 2 && DrawX == X_Pos + 14) pixel <=12'h4ff;
if (DrawY == Y_Pos + 2 && DrawX == X_Pos + 15) pixel <=12'h4ff;
if (DrawY == Y_Pos + 3 && DrawX == X_Pos + 0) pixel <=12'h4ff;
if (DrawY == Y_Pos + 3 && DrawX == X_Pos + 1) pixel <=12'h4ff;
if (DrawY == Y_Pos + 3 && DrawX == X_Pos + 2) pixel <= 12'h73f;
if (DrawY == Y_Pos + 3 && DrawX == X_Pos + 3) pixel <= 12'h73f;
if (DrawY == Y_Pos + 3 && DrawX == X_Pos + 4) pixel <= 12'h97d;
if (DrawY == Y_Pos + 3 && DrawX == X_Pos + 5) pixel <= 12'h335;
if (DrawY == Y_Pos + 3 && DrawX == X_Pos + 6) pixel <= 12'h335;
if (DrawY == Y_Pos + 3 && DrawX == X_Pos + 7) pixel <= 12'h335;
if (DrawY == Y_Pos + 3 && DrawX == X_Pos + 8) pixel <= 12'h335;
if (DrawY == Y_Pos + 3 && DrawX == X_Pos + 9) pixel <= 12'h97d;
if (DrawY == Y_Pos + 3 && DrawX == X_Pos + 10) pixel <= 12'h97d;
if (DrawY == Y_Pos + 3 && DrawX == X_Pos + 11) pixel <= 12'h73f;
if (DrawY == Y_Pos + 3 && DrawX == X_Pos + 12) pixel <= 12'h97d;
if (DrawY == Y_Pos + 3 && DrawX == X_Pos + 13) pixel <= 12'h73f;
if (DrawY == Y_Pos + 3 && DrawX == X_Pos + 14) pixel <=12'h4ff;
if (DrawY == Y_Pos + 3 && DrawX == X_Pos + 15) pixel <= 12'h73f;
if (DrawY == Y_Pos + 4 && DrawX == X_Pos + 0) pixel <=12'h4ff;
if (DrawY == Y_Pos + 4 && DrawX == X_Pos + 1) pixel <= 12'h73f;
if (DrawY == Y_Pos + 4 && DrawX == X_Pos + 2) pixel <= 12'h97d;
if (DrawY == Y_Pos + 4 && DrawX == X_Pos + 3) pixel <= 12'h335;
if (DrawY == Y_Pos + 4 && DrawX == X_Pos + 4) pixel <= 12'h335;
if (DrawY == Y_Pos + 4 && DrawX == X_Pos + 5) pixel <= 12'h335;
if (DrawY == Y_Pos + 4 && DrawX == X_Pos + 6) pixel <= 12'h335;
if (DrawY == Y_Pos + 4 && DrawX == X_Pos + 7) pixel <= 12'h224;
if (DrawY == Y_Pos + 4 && DrawX == X_Pos + 8) pixel <= 12'h224;
if (DrawY == Y_Pos + 4 && DrawX == X_Pos + 9) pixel <= 12'h224;
if (DrawY == Y_Pos + 4 && DrawX == X_Pos + 10) pixel <= 12'h224;
if (DrawY == Y_Pos + 4 && DrawX == X_Pos + 11) pixel <= 12'h97d;
if (DrawY == Y_Pos + 4 && DrawX == X_Pos + 12) pixel <=12'h4ff;
if (DrawY == Y_Pos + 4 && DrawX == X_Pos + 13) pixel <= 12'h73f;
if (DrawY == Y_Pos + 4 && DrawX == X_Pos + 14) pixel <=12'h4ff;
if (DrawY == Y_Pos + 4 && DrawX == X_Pos + 15) pixel <=12'h4ff;
if (DrawY == Y_Pos + 5 && DrawX == X_Pos + 0) pixel <=12'h4ff;
if (DrawY == Y_Pos + 5 && DrawX == X_Pos + 1) pixel <= 12'h73f;
if (DrawY == Y_Pos + 5 && DrawX == X_Pos + 2) pixel <= 12'hFFF;
if (DrawY == Y_Pos + 5 && DrawX == X_Pos + 3) pixel <= 12'h335;
if (DrawY == Y_Pos + 5 && DrawX == X_Pos + 4) pixel <= 12'h224;
if (DrawY == Y_Pos + 5 && DrawX == X_Pos + 5) pixel <= 12'h224;
if (DrawY == Y_Pos + 5 && DrawX == X_Pos + 6) pixel <= 12'h224;
if (DrawY == Y_Pos + 5 && DrawX == X_Pos + 7) pixel <= 12'h224;
if (DrawY == Y_Pos + 5 && DrawX == X_Pos + 8) pixel <= 12'h224;
if (DrawY == Y_Pos + 5 && DrawX == X_Pos + 9) pixel <= 12'h224;
if (DrawY == Y_Pos + 5 && DrawX == X_Pos + 10) pixel <= 12'h224;
if (DrawY == Y_Pos + 5 && DrawX == X_Pos + 11) pixel <= 12'hFFF;
if (DrawY == Y_Pos + 5 && DrawX == X_Pos + 12) pixel <= 12'h97d;
if (DrawY == Y_Pos + 5 && DrawX == X_Pos + 13) pixel <= 12'h73f;
if (DrawY == Y_Pos + 5 && DrawX == X_Pos + 14) pixel <= 12'h73f;
if (DrawY == Y_Pos + 5 && DrawX == X_Pos + 15) pixel <=12'h4ff;
if (DrawY == Y_Pos + 6 && DrawX == X_Pos + 0) pixel <= 12'h73f;
if (DrawY == Y_Pos + 6 && DrawX == X_Pos + 1) pixel <= 12'hFFF;
if (DrawY == Y_Pos + 6 && DrawX == X_Pos + 2) pixel <= 12'hFFF;
if (DrawY == Y_Pos + 6 && DrawX == X_Pos + 3) pixel <= 12'h335;
if (DrawY == Y_Pos + 6 && DrawX == X_Pos + 4) pixel <= 12'h224;
if (DrawY == Y_Pos + 6 && DrawX == X_Pos + 5) pixel <= 12'h224;
if (DrawY == Y_Pos + 6 && DrawX == X_Pos + 6) pixel <= 12'h224;
if (DrawY == Y_Pos + 6 && DrawX == X_Pos + 7) pixel <= 12'h224;
if (DrawY == Y_Pos + 6 && DrawX == X_Pos + 8) pixel <= 12'h224;
if (DrawY == Y_Pos + 6 && DrawX == X_Pos + 9) pixel <= 12'h224;
if (DrawY == Y_Pos + 6 && DrawX == X_Pos + 10) pixel <= 12'hFFF;
if (DrawY == Y_Pos + 6 && DrawX == X_Pos + 11) pixel <= 12'hFFF;
if (DrawY == Y_Pos + 6 && DrawX == X_Pos + 12) pixel <= 12'h224;
if (DrawY == Y_Pos + 6 && DrawX == X_Pos + 13) pixel <= 12'h97d;
if (DrawY == Y_Pos + 6 && DrawX == X_Pos + 14) pixel <=12'h4ff;
if (DrawY == Y_Pos + 6 && DrawX == X_Pos + 15) pixel <=12'h4ff;
if (DrawY == Y_Pos + 7 && DrawX == X_Pos + 0) pixel <=12'h4ff;
if (DrawY == Y_Pos + 7 && DrawX == X_Pos + 1) pixel <= 12'hFFF;
if (DrawY == Y_Pos + 7 && DrawX == X_Pos + 2) pixel <= 12'hFFF;
if (DrawY == Y_Pos + 7 && DrawX == X_Pos + 3) pixel <= 12'hFFF;
if (DrawY == Y_Pos + 7 && DrawX == X_Pos + 4) pixel <= 12'h224;
if (DrawY == Y_Pos + 7 && DrawX == X_Pos + 5) pixel <= 12'h224;
if (DrawY == Y_Pos + 7 && DrawX == X_Pos + 6) pixel <= 12'h224;
if (DrawY == Y_Pos + 7 && DrawX == X_Pos + 7) pixel <= 12'h224;
if (DrawY == Y_Pos + 7 && DrawX == X_Pos + 8) pixel <= 12'hFFF;
if (DrawY == Y_Pos + 7 && DrawX == X_Pos + 9) pixel <= 12'hFFF;
if (DrawY == Y_Pos + 7 && DrawX == X_Pos + 10) pixel <= 12'hFFF;
if (DrawY == Y_Pos + 7 && DrawX == X_Pos + 11) pixel <= 12'hFFF;
if (DrawY == Y_Pos + 7 && DrawX == X_Pos + 12) pixel <= 12'h224;
if (DrawY == Y_Pos + 7 && DrawX == X_Pos + 13) pixel <= 12'h97d;
if (DrawY == Y_Pos + 7 && DrawX == X_Pos + 14) pixel <= 12'h73f;
if (DrawY == Y_Pos + 7 && DrawX == X_Pos + 15) pixel <=12'h4ff;
if (DrawY == Y_Pos + 8 && DrawX == X_Pos + 0) pixel <=12'h4ff;
if (DrawY == Y_Pos + 8 && DrawX == X_Pos + 1) pixel <= 12'hFFF;
if (DrawY == Y_Pos + 8 && DrawX == X_Pos + 2) pixel <=12'h000;
if (DrawY == Y_Pos + 8 && DrawX == X_Pos + 3) pixel <= 12'hFFF;
if (DrawY == Y_Pos + 8 && DrawX == X_Pos + 4) pixel <= 12'hFFF;
if (DrawY == Y_Pos + 8 && DrawX == X_Pos + 5) pixel <= 12'h224;
if (DrawY == Y_Pos + 8 && DrawX == X_Pos + 6) pixel <= 12'h224;
if (DrawY == Y_Pos + 8 && DrawX == X_Pos + 7) pixel <= 12'hFFF;
if (DrawY == Y_Pos + 8 && DrawX == X_Pos + 8) pixel <=12'h000;
if (DrawY == Y_Pos + 8 && DrawX == X_Pos + 9) pixel <= 12'hFFF;
if (DrawY == Y_Pos + 8 && DrawX == X_Pos + 10) pixel <= 12'hFFF;
if (DrawY == Y_Pos + 8 && DrawX == X_Pos + 11) pixel <= 12'h224;
if (DrawY == Y_Pos + 8 && DrawX == X_Pos + 12) pixel <= 12'h224;
if (DrawY == Y_Pos + 8 && DrawX == X_Pos + 13) pixel <= 12'h97d;
if (DrawY == Y_Pos + 8 && DrawX == X_Pos + 14) pixel <= 12'h73f;
if (DrawY == Y_Pos + 8 && DrawX == X_Pos + 15) pixel <=12'h4ff;
if (DrawY == Y_Pos + 9 && DrawX == X_Pos + 0) pixel <=12'h4ff;
if (DrawY == Y_Pos + 9 && DrawX == X_Pos + 1) pixel <= 12'h73f;
if (DrawY == Y_Pos + 9 && DrawX == X_Pos + 2) pixel <= 12'hFFF;
if (DrawY == Y_Pos + 9 && DrawX == X_Pos + 3) pixel <= 12'hFFF;
if (DrawY == Y_Pos + 9 && DrawX == X_Pos + 4) pixel <= 12'h224;
if (DrawY == Y_Pos + 9 && DrawX == X_Pos + 5) pixel <= 12'h224;
if (DrawY == Y_Pos + 9 && DrawX == X_Pos + 6) pixel <= 12'h224;
if (DrawY == Y_Pos + 9 && DrawX == X_Pos + 7) pixel <= 12'h224;
if (DrawY == Y_Pos + 9 && DrawX == X_Pos + 8) pixel <= 12'hFFF;
if (DrawY == Y_Pos + 9 && DrawX == X_Pos + 9) pixel <= 12'hFFF;
if (DrawY == Y_Pos + 9 && DrawX == X_Pos + 10) pixel <= 12'h224;
if (DrawY == Y_Pos + 9 && DrawX == X_Pos + 11) pixel <= 12'h224;
if (DrawY == Y_Pos + 9 && DrawX == X_Pos + 12) pixel <= 12'h224;
if (DrawY == Y_Pos + 9 && DrawX == X_Pos + 13) pixel <= 12'h97d;
if (DrawY == Y_Pos + 9 && DrawX == X_Pos + 14) pixel <= 12'h73f;
if (DrawY == Y_Pos + 9 && DrawX == X_Pos + 15) pixel <=12'h4ff;
if (DrawY == Y_Pos + 10 && DrawX == X_Pos + 0) pixel <= 12'h73f;
if (DrawY == Y_Pos + 10 && DrawX == X_Pos + 1) pixel <= 12'h73f;
if (DrawY == Y_Pos + 10 && DrawX == X_Pos + 2) pixel <= 12'h224;
if (DrawY == Y_Pos + 10 && DrawX == X_Pos + 3) pixel <= 12'h224;
if (DrawY == Y_Pos + 10 && DrawX == X_Pos + 4) pixel <= 12'h224;
if (DrawY == Y_Pos + 10 && DrawX == X_Pos + 5) pixel <= 12'h224;
if (DrawY == Y_Pos + 10 && DrawX == X_Pos + 6) pixel <= 12'h224;
if (DrawY == Y_Pos + 10 && DrawX == X_Pos + 7) pixel <= 12'h224;
if (DrawY == Y_Pos + 10 && DrawX == X_Pos + 8) pixel <= 12'h224;
if (DrawY == Y_Pos + 10 && DrawX == X_Pos + 9) pixel <= 12'h224;
if (DrawY == Y_Pos + 10 && DrawX == X_Pos + 10) pixel <= 12'h224;
if (DrawY == Y_Pos + 10 && DrawX == X_Pos + 11) pixel <= 12'h224;
if (DrawY == Y_Pos + 10 && DrawX == X_Pos + 12) pixel <= 12'h224;
if (DrawY == Y_Pos + 10 && DrawX == X_Pos + 13) pixel <= 12'h97d;
if (DrawY == Y_Pos + 10 && DrawX == X_Pos + 14) pixel <=12'h4ff;
if (DrawY == Y_Pos + 10 && DrawX == X_Pos + 15) pixel <= 12'h73f;
if (DrawY == Y_Pos + 11 && DrawX == X_Pos + 0) pixel <=12'h4ff;
if (DrawY == Y_Pos + 11 && DrawX == X_Pos + 1) pixel <= 12'h73f;
if (DrawY == Y_Pos + 11 && DrawX == X_Pos + 2) pixel <= 12'h73f;
if (DrawY == Y_Pos + 11 && DrawX == X_Pos + 3) pixel <= 12'hFFF;
if (DrawY == Y_Pos + 11 && DrawX == X_Pos + 4) pixel <= 12'hd79;
if (DrawY == Y_Pos + 11 && DrawX == X_Pos + 5) pixel <= 12'hd79;
if (DrawY == Y_Pos + 11 && DrawX == X_Pos + 6) pixel <= 12'hd79;
if (DrawY == Y_Pos + 11 && DrawX == X_Pos + 7) pixel <= 12'hd79;
if (DrawY == Y_Pos + 11 && DrawX == X_Pos + 8) pixel <= 12'hFFF;
if (DrawY == Y_Pos + 11 && DrawX == X_Pos + 9) pixel <= 12'h224;
if (DrawY == Y_Pos + 11 && DrawX == X_Pos + 10) pixel <= 12'h224;
if (DrawY == Y_Pos + 11 && DrawX == X_Pos + 11) pixel <= 12'h224;
if (DrawY == Y_Pos + 11 && DrawX == X_Pos + 12) pixel <= 12'h97d;
if (DrawY == Y_Pos + 11 && DrawX == X_Pos + 13) pixel <= 12'h73f;
if (DrawY == Y_Pos + 11 && DrawX == X_Pos + 14) pixel <=12'h4ff;
if (DrawY == Y_Pos + 11 && DrawX == X_Pos + 15) pixel <=12'h4ff;
if (DrawY == Y_Pos + 12 && DrawX == X_Pos + 0) pixel <=12'h4ff;
if (DrawY == Y_Pos + 12 && DrawX == X_Pos + 1) pixel <=12'h4ff;
if (DrawY == Y_Pos + 12 && DrawX == X_Pos + 2) pixel <= 12'h73f;
if (DrawY == Y_Pos + 12 && DrawX == X_Pos + 3) pixel <= 12'hFFF;
if (DrawY == Y_Pos + 12 && DrawX == X_Pos + 4) pixel <= 12'h335;
if (DrawY == Y_Pos + 12 && DrawX == X_Pos + 5) pixel <= 12'h335;
if (DrawY == Y_Pos + 12 && DrawX == X_Pos + 6) pixel <= 12'h224;
if (DrawY == Y_Pos + 12 && DrawX == X_Pos + 7) pixel <= 12'h224;
if (DrawY == Y_Pos + 12 && DrawX == X_Pos + 8) pixel <= 12'hFFF;
if (DrawY == Y_Pos + 12 && DrawX == X_Pos + 9) pixel <= 12'h224;
if (DrawY == Y_Pos + 12 && DrawX == X_Pos + 10) pixel <= 12'h224;
if (DrawY == Y_Pos + 12 && DrawX == X_Pos + 11) pixel <= 12'h97d;
if (DrawY == Y_Pos + 12 && DrawX == X_Pos + 12) pixel <= 12'h73f;
if (DrawY == Y_Pos + 12 && DrawX == X_Pos + 13) pixel <=12'h4ff;
if (DrawY == Y_Pos + 12 && DrawX == X_Pos + 14) pixel <=12'h4ff;
if (DrawY == Y_Pos + 12 && DrawX == X_Pos + 15) pixel <=12'h4ff;
if (DrawY == Y_Pos + 13 && DrawX == X_Pos + 0) pixel <=12'h4ff;
if (DrawY == Y_Pos + 13 && DrawX == X_Pos + 1) pixel <=12'h4ff;
if (DrawY == Y_Pos + 13 && DrawX == X_Pos + 2) pixel <=12'h4ff;
if (DrawY == Y_Pos + 13 && DrawX == X_Pos + 3) pixel <= 12'h73f;
if (DrawY == Y_Pos + 13 && DrawX == X_Pos + 4) pixel <= 12'h73f;
if (DrawY == Y_Pos + 13 && DrawX == X_Pos + 5) pixel <= 12'h335;
if (DrawY == Y_Pos + 13 && DrawX == X_Pos + 6) pixel <= 12'h335;
if (DrawY == Y_Pos + 13 && DrawX == X_Pos + 7) pixel <= 12'h335;
if (DrawY == Y_Pos + 13 && DrawX == X_Pos + 8) pixel <= 12'h224;
if (DrawY == Y_Pos + 13 && DrawX == X_Pos + 9) pixel <= 12'h97d;
if (DrawY == Y_Pos + 13 && DrawX == X_Pos + 10) pixel <= 12'h73f;
if (DrawY == Y_Pos + 13 && DrawX == X_Pos + 11) pixel <=12'h4ff;
if (DrawY == Y_Pos + 13 && DrawX == X_Pos + 12) pixel <=12'h4ff;
if (DrawY == Y_Pos + 13 && DrawX == X_Pos + 13) pixel <= 12'h73f;
if (DrawY == Y_Pos + 13 && DrawX == X_Pos + 14) pixel <= 12'h73f;
if (DrawY == Y_Pos + 13 && DrawX == X_Pos + 15) pixel <=12'h4ff;
if (DrawY == Y_Pos + 14 && DrawX == X_Pos + 0) pixel <=12'h4ff;
if (DrawY == Y_Pos + 14 && DrawX == X_Pos + 1) pixel <=12'h4ff;
if (DrawY == Y_Pos + 14 && DrawX == X_Pos + 2) pixel <= 12'h73f;
if (DrawY == Y_Pos + 14 && DrawX == X_Pos + 3) pixel <=12'h4ff;
if (DrawY == Y_Pos + 14 && DrawX == X_Pos + 4) pixel <=12'h4ff;
if (DrawY == Y_Pos + 14 && DrawX == X_Pos + 5) pixel <= 12'h73f;
if (DrawY == Y_Pos + 14 && DrawX == X_Pos + 6) pixel <= 12'h73f;
if (DrawY == Y_Pos + 14 && DrawX == X_Pos + 7) pixel <= 12'h97d;
if (DrawY == Y_Pos + 14 && DrawX == X_Pos + 8) pixel <= 12'h97d;
if (DrawY == Y_Pos + 14 && DrawX == X_Pos + 9) pixel <= 12'h73f;
if (DrawY == Y_Pos + 14 && DrawX == X_Pos + 10) pixel <= 12'h73f;
if (DrawY == Y_Pos + 14 && DrawX == X_Pos + 11) pixel <=12'h4ff;
if (DrawY == Y_Pos + 14 && DrawX == X_Pos + 12) pixel <=12'h4ff;
if (DrawY == Y_Pos + 14 && DrawX == X_Pos + 13) pixel <=12'h4ff;
if (DrawY == Y_Pos + 14 && DrawX == X_Pos + 14) pixel <=12'h4ff;
if (DrawY == Y_Pos + 14 && DrawX == X_Pos + 15) pixel <= 12'h73f;
if (DrawY == Y_Pos + 15 && DrawX == X_Pos + 0) pixel <=12'h4ff;
if (DrawY == Y_Pos + 15 && DrawX == X_Pos + 1) pixel <=12'h4ff;
if (DrawY == Y_Pos + 15 && DrawX == X_Pos + 2) pixel <=12'h4ff;
if (DrawY == Y_Pos + 15 && DrawX == X_Pos + 3) pixel <=12'h4ff;
if (DrawY == Y_Pos + 15 && DrawX == X_Pos + 4) pixel <=12'h4ff;
if (DrawY == Y_Pos + 15 && DrawX == X_Pos + 5) pixel <=12'h4ff;
if (DrawY == Y_Pos + 15 && DrawX == X_Pos + 6) pixel <=12'h4ff;
if (DrawY == Y_Pos + 15 && DrawX == X_Pos + 7) pixel <= 12'h73f;
if (DrawY == Y_Pos + 15 && DrawX == X_Pos + 8) pixel <=12'h4ff;
if (DrawY == Y_Pos + 15 && DrawX == X_Pos + 9) pixel <=12'h4ff;
if (DrawY == Y_Pos + 15 && DrawX == X_Pos + 10) pixel <=12'h4ff;
if (DrawY == Y_Pos + 15 && DrawX == X_Pos + 11) pixel <= 12'h73f;
if (DrawY == Y_Pos + 15 && DrawX == X_Pos + 12) pixel <=12'h4ff;
if (DrawY == Y_Pos + 15 && DrawX == X_Pos + 13) pixel <=12'h4ff;
if (DrawY == Y_Pos + 15 && DrawX == X_Pos + 14) pixel <=12'h4ff;
if (DrawY == Y_Pos + 15 && DrawX == X_Pos + 15) pixel <=12'h4ff;
else pixel <=12'h4ff;