module pacman_wall_collision (
	input logic [9:0] X_Pos,
	input logic [9:0] Y_Pos,

	output logic Is_Wall);

always_comb begin
	Is_Wall = 1'b0;

	if ((X_Pos > 10'd125) && (X_Pos < 10'd514) && (Y_Pos > 10'd46) && (Y_Pos < 10'd50)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd125) && (X_Pos < 10'd514) && (Y_Pos > 10'd47) && (Y_Pos < 10'd51)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd122) && (X_Pos < 10'd128) && (Y_Pos > 10'd48) && (Y_Pos < 10'd52)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd517) && (Y_Pos > 10'd48) && (Y_Pos < 10'd52)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd120) && (X_Pos < 10'd125) && (Y_Pos > 10'd49) && (Y_Pos < 10'd53)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd514) && (X_Pos < 10'd519) && (Y_Pos > 10'd49) && (Y_Pos < 10'd53)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd120) && (X_Pos < 10'd125) && (Y_Pos > 10'd50) && (Y_Pos < 10'd54)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd514) && (X_Pos < 10'd519) && (Y_Pos > 10'd50) && (Y_Pos < 10'd54)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd120) && (X_Pos < 10'd125) && (Y_Pos > 10'd51) && (Y_Pos < 10'd55)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd127) && (X_Pos < 10'd312) && (Y_Pos > 10'd51) && (Y_Pos < 10'd55)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd327) && (X_Pos < 10'd512) && (Y_Pos > 10'd51) && (Y_Pos < 10'd55)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd514) && (X_Pos < 10'd519) && (Y_Pos > 10'd51) && (Y_Pos < 10'd55)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd52) && (Y_Pos < 10'd56)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd125) && (X_Pos < 10'd314) && (Y_Pos > 10'd52) && (Y_Pos < 10'd56)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd325) && (X_Pos < 10'd514) && (Y_Pos > 10'd52) && (Y_Pos < 10'd56)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd52) && (Y_Pos < 10'd56)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd53) && (Y_Pos < 10'd57)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd125) && (X_Pos < 10'd130) && (Y_Pos > 10'd53) && (Y_Pos < 10'd57)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd309) && (X_Pos < 10'd314) && (Y_Pos > 10'd53) && (Y_Pos < 10'd57)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd325) && (X_Pos < 10'd330) && (Y_Pos > 10'd53) && (Y_Pos < 10'd57)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd509) && (X_Pos < 10'd514) && (Y_Pos > 10'd53) && (Y_Pos < 10'd57)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd53) && (Y_Pos < 10'd57)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd54) && (Y_Pos < 10'd58)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd54) && (Y_Pos < 10'd58)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd54) && (Y_Pos < 10'd58)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd54) && (Y_Pos < 10'd58)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd54) && (Y_Pos < 10'd58)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd54) && (Y_Pos < 10'd58)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd55) && (Y_Pos < 10'd59)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd55) && (Y_Pos < 10'd59)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd55) && (Y_Pos < 10'd59)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd55) && (Y_Pos < 10'd59)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd55) && (Y_Pos < 10'd59)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd55) && (Y_Pos < 10'd59)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd56) && (Y_Pos < 10'd60)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd56) && (Y_Pos < 10'd60)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd56) && (Y_Pos < 10'd60)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd56) && (Y_Pos < 10'd60)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd56) && (Y_Pos < 10'd60)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd56) && (Y_Pos < 10'd60)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd57) && (Y_Pos < 10'd61)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd57) && (Y_Pos < 10'd61)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd57) && (Y_Pos < 10'd61)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd57) && (Y_Pos < 10'd61)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd57) && (Y_Pos < 10'd61)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd57) && (Y_Pos < 10'd61)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd58) && (Y_Pos < 10'd62)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd58) && (Y_Pos < 10'd62)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd58) && (Y_Pos < 10'd62)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd58) && (Y_Pos < 10'd62)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd58) && (Y_Pos < 10'd62)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd58) && (Y_Pos < 10'd62)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd59) && (Y_Pos < 10'd63)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd59) && (Y_Pos < 10'd63)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd59) && (Y_Pos < 10'd63)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd59) && (Y_Pos < 10'd63)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd59) && (Y_Pos < 10'd63)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd59) && (Y_Pos < 10'd63)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd60) && (Y_Pos < 10'd64)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd60) && (Y_Pos < 10'd64)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd60) && (Y_Pos < 10'd64)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd60) && (Y_Pos < 10'd64)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd60) && (Y_Pos < 10'd64)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd60) && (Y_Pos < 10'd64)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd61) && (Y_Pos < 10'd65)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd61) && (Y_Pos < 10'd65)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd61) && (Y_Pos < 10'd65)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd61) && (Y_Pos < 10'd65)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd61) && (Y_Pos < 10'd65)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd61) && (Y_Pos < 10'd65)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd62) && (Y_Pos < 10'd66)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd62) && (Y_Pos < 10'd66)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd62) && (Y_Pos < 10'd66)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd62) && (Y_Pos < 10'd66)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd62) && (Y_Pos < 10'd66)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd62) && (Y_Pos < 10'd66)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd63) && (Y_Pos < 10'd67)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd63) && (Y_Pos < 10'd67)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd63) && (Y_Pos < 10'd67)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd63) && (Y_Pos < 10'd67)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd63) && (Y_Pos < 10'd67)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd63) && (Y_Pos < 10'd67)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd64) && (Y_Pos < 10'd68)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd64) && (Y_Pos < 10'd68)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd64) && (Y_Pos < 10'd68)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd64) && (Y_Pos < 10'd68)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd64) && (Y_Pos < 10'd68)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd64) && (Y_Pos < 10'd68)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd65) && (Y_Pos < 10'd69)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd65) && (Y_Pos < 10'd69)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd65) && (Y_Pos < 10'd69)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd65) && (Y_Pos < 10'd69)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd65) && (Y_Pos < 10'd69)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd65) && (Y_Pos < 10'd69)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd66) && (Y_Pos < 10'd70)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd66) && (Y_Pos < 10'd70)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd66) && (Y_Pos < 10'd70)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd66) && (Y_Pos < 10'd70)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd66) && (Y_Pos < 10'd70)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd66) && (Y_Pos < 10'd70)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd67) && (Y_Pos < 10'd71)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd67) && (Y_Pos < 10'd71)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd67) && (Y_Pos < 10'd71)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd67) && (Y_Pos < 10'd71)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd67) && (Y_Pos < 10'd71)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd67) && (Y_Pos < 10'd71)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd68) && (Y_Pos < 10'd72)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd68) && (Y_Pos < 10'd72)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd68) && (Y_Pos < 10'd72)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd68) && (Y_Pos < 10'd72)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd68) && (Y_Pos < 10'd72)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd68) && (Y_Pos < 10'd72)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd69) && (Y_Pos < 10'd73)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd69) && (Y_Pos < 10'd73)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd69) && (Y_Pos < 10'd73)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd69) && (Y_Pos < 10'd73)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd69) && (Y_Pos < 10'd73)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd69) && (Y_Pos < 10'd73)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd70) && (Y_Pos < 10'd74)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd70) && (Y_Pos < 10'd74)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd70) && (Y_Pos < 10'd74)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd70) && (Y_Pos < 10'd74)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd70) && (Y_Pos < 10'd74)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd70) && (Y_Pos < 10'd74)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd71) && (Y_Pos < 10'd75)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd71) && (Y_Pos < 10'd75)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd71) && (Y_Pos < 10'd75)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd71) && (Y_Pos < 10'd75)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd71) && (Y_Pos < 10'd75)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd71) && (Y_Pos < 10'd75)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd72) && (Y_Pos < 10'd76)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd72) && (Y_Pos < 10'd76)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd72) && (Y_Pos < 10'd76)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd72) && (Y_Pos < 10'd76)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd72) && (Y_Pos < 10'd76)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd72) && (Y_Pos < 10'd76)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd73) && (Y_Pos < 10'd77)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd73) && (Y_Pos < 10'd77)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd73) && (Y_Pos < 10'd77)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd73) && (Y_Pos < 10'd77)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd73) && (Y_Pos < 10'd77)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd73) && (Y_Pos < 10'd77)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd74) && (Y_Pos < 10'd78)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd74) && (Y_Pos < 10'd78)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd74) && (Y_Pos < 10'd78)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd74) && (Y_Pos < 10'd78)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd74) && (Y_Pos < 10'd78)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd74) && (Y_Pos < 10'd78)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd75) && (Y_Pos < 10'd79)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd75) && (Y_Pos < 10'd79)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd75) && (Y_Pos < 10'd79)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd75) && (Y_Pos < 10'd79)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd75) && (Y_Pos < 10'd79)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd75) && (Y_Pos < 10'd79)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd76) && (Y_Pos < 10'd80)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd76) && (Y_Pos < 10'd80)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd76) && (Y_Pos < 10'd80)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd76) && (Y_Pos < 10'd80)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd76) && (Y_Pos < 10'd80)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd76) && (Y_Pos < 10'd80)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd77) && (Y_Pos < 10'd81)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd77) && (Y_Pos < 10'd81)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd77) && (Y_Pos < 10'd81)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd77) && (Y_Pos < 10'd81)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd77) && (Y_Pos < 10'd81)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd77) && (Y_Pos < 10'd81)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd78) && (Y_Pos < 10'd82)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd78) && (Y_Pos < 10'd82)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd158) && (X_Pos < 10'd196) && (Y_Pos > 10'd78) && (Y_Pos < 10'd82)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd229) && (X_Pos < 10'd281) && (Y_Pos > 10'd78) && (Y_Pos < 10'd82)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd78) && (Y_Pos < 10'd82)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd78) && (Y_Pos < 10'd82)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd358) && (X_Pos < 10'd410) && (Y_Pos > 10'd78) && (Y_Pos < 10'd82)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd443) && (X_Pos < 10'd481) && (Y_Pos > 10'd78) && (Y_Pos < 10'd82)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd78) && (Y_Pos < 10'd82)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd78) && (Y_Pos < 10'd82)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd79) && (Y_Pos < 10'd83)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd79) && (Y_Pos < 10'd83)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd157) && (X_Pos < 10'd196) && (Y_Pos > 10'd79) && (Y_Pos < 10'd83)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd228) && (X_Pos < 10'd282) && (Y_Pos > 10'd79) && (Y_Pos < 10'd83)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd79) && (Y_Pos < 10'd83)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd79) && (Y_Pos < 10'd83)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd357) && (X_Pos < 10'd411) && (Y_Pos > 10'd79) && (Y_Pos < 10'd83)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd443) && (X_Pos < 10'd482) && (Y_Pos > 10'd79) && (Y_Pos < 10'd83)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd79) && (Y_Pos < 10'd83)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd79) && (Y_Pos < 10'd83)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd80) && (Y_Pos < 10'd84)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd80) && (Y_Pos < 10'd84)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd155) && (X_Pos < 10'd160) && (Y_Pos > 10'd80) && (Y_Pos < 10'd84)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd193) && (X_Pos < 10'd198) && (Y_Pos > 10'd80) && (Y_Pos < 10'd84)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd227) && (X_Pos < 10'd232) && (Y_Pos > 10'd80) && (Y_Pos < 10'd84)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd279) && (X_Pos < 10'd284) && (Y_Pos > 10'd80) && (Y_Pos < 10'd84)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd80) && (Y_Pos < 10'd84)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd80) && (Y_Pos < 10'd84)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd355) && (X_Pos < 10'd360) && (Y_Pos > 10'd80) && (Y_Pos < 10'd84)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd407) && (X_Pos < 10'd412) && (Y_Pos > 10'd80) && (Y_Pos < 10'd84)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd441) && (X_Pos < 10'd446) && (Y_Pos > 10'd80) && (Y_Pos < 10'd84)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd479) && (X_Pos < 10'd484) && (Y_Pos > 10'd80) && (Y_Pos < 10'd84)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd80) && (Y_Pos < 10'd84)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd80) && (Y_Pos < 10'd84)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd81) && (Y_Pos < 10'd85)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd81) && (Y_Pos < 10'd85)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd155) && (X_Pos < 10'd160) && (Y_Pos > 10'd81) && (Y_Pos < 10'd85)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd193) && (X_Pos < 10'd199) && (Y_Pos > 10'd81) && (Y_Pos < 10'd85)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd226) && (X_Pos < 10'd231) && (Y_Pos > 10'd81) && (Y_Pos < 10'd85)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd279) && (X_Pos < 10'd284) && (Y_Pos > 10'd81) && (Y_Pos < 10'd85)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd81) && (Y_Pos < 10'd85)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd81) && (Y_Pos < 10'd85)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd355) && (X_Pos < 10'd360) && (Y_Pos > 10'd81) && (Y_Pos < 10'd85)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd408) && (X_Pos < 10'd413) && (Y_Pos > 10'd81) && (Y_Pos < 10'd85)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd440) && (X_Pos < 10'd446) && (Y_Pos > 10'd81) && (Y_Pos < 10'd85)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd479) && (X_Pos < 10'd484) && (Y_Pos > 10'd81) && (Y_Pos < 10'd85)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd81) && (Y_Pos < 10'd85)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd81) && (Y_Pos < 10'd85)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd82) && (Y_Pos < 10'd86)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd82) && (Y_Pos < 10'd86)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd154) && (X_Pos < 10'd159) && (Y_Pos > 10'd82) && (Y_Pos < 10'd86)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd82) && (Y_Pos < 10'd86)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd82) && (Y_Pos < 10'd86)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd280) && (X_Pos < 10'd285) && (Y_Pos > 10'd82) && (Y_Pos < 10'd86)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd82) && (Y_Pos < 10'd86)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd82) && (Y_Pos < 10'd86)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd354) && (X_Pos < 10'd359) && (Y_Pos > 10'd82) && (Y_Pos < 10'd86)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd82) && (Y_Pos < 10'd86)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd82) && (Y_Pos < 10'd86)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd480) && (X_Pos < 10'd485) && (Y_Pos > 10'd82) && (Y_Pos < 10'd86)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd82) && (Y_Pos < 10'd86)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd82) && (Y_Pos < 10'd86)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd83) && (Y_Pos < 10'd87)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd83) && (Y_Pos < 10'd87)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd154) && (X_Pos < 10'd159) && (Y_Pos > 10'd83) && (Y_Pos < 10'd87)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd83) && (Y_Pos < 10'd87)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd83) && (Y_Pos < 10'd87)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd280) && (X_Pos < 10'd285) && (Y_Pos > 10'd83) && (Y_Pos < 10'd87)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd83) && (Y_Pos < 10'd87)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd83) && (Y_Pos < 10'd87)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd354) && (X_Pos < 10'd359) && (Y_Pos > 10'd83) && (Y_Pos < 10'd87)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd83) && (Y_Pos < 10'd87)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd83) && (Y_Pos < 10'd87)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd480) && (X_Pos < 10'd485) && (Y_Pos > 10'd83) && (Y_Pos < 10'd87)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd83) && (Y_Pos < 10'd87)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd83) && (Y_Pos < 10'd87)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd84) && (Y_Pos < 10'd88)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd84) && (Y_Pos < 10'd88)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd154) && (X_Pos < 10'd159) && (Y_Pos > 10'd84) && (Y_Pos < 10'd88)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd84) && (Y_Pos < 10'd88)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd84) && (Y_Pos < 10'd88)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd280) && (X_Pos < 10'd285) && (Y_Pos > 10'd84) && (Y_Pos < 10'd88)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd84) && (Y_Pos < 10'd88)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd84) && (Y_Pos < 10'd88)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd354) && (X_Pos < 10'd359) && (Y_Pos > 10'd84) && (Y_Pos < 10'd88)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd84) && (Y_Pos < 10'd88)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd84) && (Y_Pos < 10'd88)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd480) && (X_Pos < 10'd485) && (Y_Pos > 10'd84) && (Y_Pos < 10'd88)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd84) && (Y_Pos < 10'd88)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd84) && (Y_Pos < 10'd88)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd85) && (Y_Pos < 10'd89)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd85) && (Y_Pos < 10'd89)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd154) && (X_Pos < 10'd159) && (Y_Pos > 10'd85) && (Y_Pos < 10'd89)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd85) && (Y_Pos < 10'd89)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd85) && (Y_Pos < 10'd89)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd280) && (X_Pos < 10'd285) && (Y_Pos > 10'd85) && (Y_Pos < 10'd89)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd85) && (Y_Pos < 10'd89)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd85) && (Y_Pos < 10'd89)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd354) && (X_Pos < 10'd359) && (Y_Pos > 10'd85) && (Y_Pos < 10'd89)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd85) && (Y_Pos < 10'd89)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd85) && (Y_Pos < 10'd89)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd480) && (X_Pos < 10'd485) && (Y_Pos > 10'd85) && (Y_Pos < 10'd89)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd85) && (Y_Pos < 10'd89)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd85) && (Y_Pos < 10'd89)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd86) && (Y_Pos < 10'd90)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd86) && (Y_Pos < 10'd90)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd154) && (X_Pos < 10'd159) && (Y_Pos > 10'd86) && (Y_Pos < 10'd90)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd86) && (Y_Pos < 10'd90)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd86) && (Y_Pos < 10'd90)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd280) && (X_Pos < 10'd285) && (Y_Pos > 10'd86) && (Y_Pos < 10'd90)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd86) && (Y_Pos < 10'd90)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd86) && (Y_Pos < 10'd90)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd354) && (X_Pos < 10'd359) && (Y_Pos > 10'd86) && (Y_Pos < 10'd90)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd86) && (Y_Pos < 10'd90)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd86) && (Y_Pos < 10'd90)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd480) && (X_Pos < 10'd485) && (Y_Pos > 10'd86) && (Y_Pos < 10'd90)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd86) && (Y_Pos < 10'd90)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd86) && (Y_Pos < 10'd90)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd87) && (Y_Pos < 10'd91)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd87) && (Y_Pos < 10'd91)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd154) && (X_Pos < 10'd159) && (Y_Pos > 10'd87) && (Y_Pos < 10'd91)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd87) && (Y_Pos < 10'd91)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd87) && (Y_Pos < 10'd91)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd280) && (X_Pos < 10'd285) && (Y_Pos > 10'd87) && (Y_Pos < 10'd91)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd87) && (Y_Pos < 10'd91)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd87) && (Y_Pos < 10'd91)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd354) && (X_Pos < 10'd359) && (Y_Pos > 10'd87) && (Y_Pos < 10'd91)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd87) && (Y_Pos < 10'd91)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd87) && (Y_Pos < 10'd91)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd480) && (X_Pos < 10'd485) && (Y_Pos > 10'd87) && (Y_Pos < 10'd91)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd87) && (Y_Pos < 10'd91)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd87) && (Y_Pos < 10'd91)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd88) && (Y_Pos < 10'd92)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd88) && (Y_Pos < 10'd92)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd154) && (X_Pos < 10'd159) && (Y_Pos > 10'd88) && (Y_Pos < 10'd92)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd88) && (Y_Pos < 10'd92)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd88) && (Y_Pos < 10'd92)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd280) && (X_Pos < 10'd285) && (Y_Pos > 10'd88) && (Y_Pos < 10'd92)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd88) && (Y_Pos < 10'd92)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd88) && (Y_Pos < 10'd92)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd354) && (X_Pos < 10'd359) && (Y_Pos > 10'd88) && (Y_Pos < 10'd92)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd88) && (Y_Pos < 10'd92)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd88) && (Y_Pos < 10'd92)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd480) && (X_Pos < 10'd485) && (Y_Pos > 10'd88) && (Y_Pos < 10'd92)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd88) && (Y_Pos < 10'd92)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd88) && (Y_Pos < 10'd92)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd89) && (Y_Pos < 10'd93)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd89) && (Y_Pos < 10'd93)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd154) && (X_Pos < 10'd159) && (Y_Pos > 10'd89) && (Y_Pos < 10'd93)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd89) && (Y_Pos < 10'd93)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd89) && (Y_Pos < 10'd93)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd280) && (X_Pos < 10'd285) && (Y_Pos > 10'd89) && (Y_Pos < 10'd93)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd89) && (Y_Pos < 10'd93)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd89) && (Y_Pos < 10'd93)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd354) && (X_Pos < 10'd359) && (Y_Pos > 10'd89) && (Y_Pos < 10'd93)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd89) && (Y_Pos < 10'd93)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd89) && (Y_Pos < 10'd93)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd480) && (X_Pos < 10'd485) && (Y_Pos > 10'd89) && (Y_Pos < 10'd93)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd89) && (Y_Pos < 10'd93)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd89) && (Y_Pos < 10'd93)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd90) && (Y_Pos < 10'd94)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd90) && (Y_Pos < 10'd94)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd154) && (X_Pos < 10'd159) && (Y_Pos > 10'd90) && (Y_Pos < 10'd94)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd90) && (Y_Pos < 10'd94)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd90) && (Y_Pos < 10'd94)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd280) && (X_Pos < 10'd285) && (Y_Pos > 10'd90) && (Y_Pos < 10'd94)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd90) && (Y_Pos < 10'd94)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd90) && (Y_Pos < 10'd94)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd354) && (X_Pos < 10'd359) && (Y_Pos > 10'd90) && (Y_Pos < 10'd94)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd90) && (Y_Pos < 10'd94)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd90) && (Y_Pos < 10'd94)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd480) && (X_Pos < 10'd485) && (Y_Pos > 10'd90) && (Y_Pos < 10'd94)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd90) && (Y_Pos < 10'd94)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd90) && (Y_Pos < 10'd94)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd91) && (Y_Pos < 10'd95)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd91) && (Y_Pos < 10'd95)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd154) && (X_Pos < 10'd159) && (Y_Pos > 10'd91) && (Y_Pos < 10'd95)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd91) && (Y_Pos < 10'd95)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd91) && (Y_Pos < 10'd95)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd280) && (X_Pos < 10'd285) && (Y_Pos > 10'd91) && (Y_Pos < 10'd95)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd91) && (Y_Pos < 10'd95)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd91) && (Y_Pos < 10'd95)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd354) && (X_Pos < 10'd359) && (Y_Pos > 10'd91) && (Y_Pos < 10'd95)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd91) && (Y_Pos < 10'd95)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd91) && (Y_Pos < 10'd95)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd480) && (X_Pos < 10'd485) && (Y_Pos > 10'd91) && (Y_Pos < 10'd95)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd91) && (Y_Pos < 10'd95)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd91) && (Y_Pos < 10'd95)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd92) && (Y_Pos < 10'd96)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd92) && (Y_Pos < 10'd96)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd154) && (X_Pos < 10'd159) && (Y_Pos > 10'd92) && (Y_Pos < 10'd96)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd92) && (Y_Pos < 10'd96)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd92) && (Y_Pos < 10'd96)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd280) && (X_Pos < 10'd285) && (Y_Pos > 10'd92) && (Y_Pos < 10'd96)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd92) && (Y_Pos < 10'd96)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd92) && (Y_Pos < 10'd96)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd354) && (X_Pos < 10'd359) && (Y_Pos > 10'd92) && (Y_Pos < 10'd96)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd92) && (Y_Pos < 10'd96)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd92) && (Y_Pos < 10'd96)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd480) && (X_Pos < 10'd485) && (Y_Pos > 10'd92) && (Y_Pos < 10'd96)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd92) && (Y_Pos < 10'd96)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd92) && (Y_Pos < 10'd96)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd93) && (Y_Pos < 10'd97)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd93) && (Y_Pos < 10'd97)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd154) && (X_Pos < 10'd159) && (Y_Pos > 10'd93) && (Y_Pos < 10'd97)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd93) && (Y_Pos < 10'd97)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd93) && (Y_Pos < 10'd97)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd280) && (X_Pos < 10'd285) && (Y_Pos > 10'd93) && (Y_Pos < 10'd97)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd93) && (Y_Pos < 10'd97)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd93) && (Y_Pos < 10'd97)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd354) && (X_Pos < 10'd359) && (Y_Pos > 10'd93) && (Y_Pos < 10'd97)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd93) && (Y_Pos < 10'd97)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd93) && (Y_Pos < 10'd97)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd480) && (X_Pos < 10'd485) && (Y_Pos > 10'd93) && (Y_Pos < 10'd97)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd93) && (Y_Pos < 10'd97)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd93) && (Y_Pos < 10'd97)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd94) && (Y_Pos < 10'd98)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd94) && (Y_Pos < 10'd98)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd154) && (X_Pos < 10'd159) && (Y_Pos > 10'd94) && (Y_Pos < 10'd98)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd94) && (Y_Pos < 10'd98)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd94) && (Y_Pos < 10'd98)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd280) && (X_Pos < 10'd285) && (Y_Pos > 10'd94) && (Y_Pos < 10'd98)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd94) && (Y_Pos < 10'd98)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd94) && (Y_Pos < 10'd98)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd354) && (X_Pos < 10'd359) && (Y_Pos > 10'd94) && (Y_Pos < 10'd98)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd94) && (Y_Pos < 10'd98)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd94) && (Y_Pos < 10'd98)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd480) && (X_Pos < 10'd485) && (Y_Pos > 10'd94) && (Y_Pos < 10'd98)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd94) && (Y_Pos < 10'd98)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd94) && (Y_Pos < 10'd98)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd95) && (Y_Pos < 10'd99)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd95) && (Y_Pos < 10'd99)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd154) && (X_Pos < 10'd159) && (Y_Pos > 10'd95) && (Y_Pos < 10'd99)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd95) && (Y_Pos < 10'd99)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd95) && (Y_Pos < 10'd99)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd280) && (X_Pos < 10'd285) && (Y_Pos > 10'd95) && (Y_Pos < 10'd99)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd95) && (Y_Pos < 10'd99)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd95) && (Y_Pos < 10'd99)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd354) && (X_Pos < 10'd359) && (Y_Pos > 10'd95) && (Y_Pos < 10'd99)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd95) && (Y_Pos < 10'd99)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd95) && (Y_Pos < 10'd99)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd480) && (X_Pos < 10'd485) && (Y_Pos > 10'd95) && (Y_Pos < 10'd99)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd95) && (Y_Pos < 10'd99)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd95) && (Y_Pos < 10'd99)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd96) && (Y_Pos < 10'd100)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd96) && (Y_Pos < 10'd100)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd154) && (X_Pos < 10'd159) && (Y_Pos > 10'd96) && (Y_Pos < 10'd100)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd96) && (Y_Pos < 10'd100)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd96) && (Y_Pos < 10'd100)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd280) && (X_Pos < 10'd285) && (Y_Pos > 10'd96) && (Y_Pos < 10'd100)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd96) && (Y_Pos < 10'd100)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd96) && (Y_Pos < 10'd100)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd354) && (X_Pos < 10'd359) && (Y_Pos > 10'd96) && (Y_Pos < 10'd100)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd96) && (Y_Pos < 10'd100)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd96) && (Y_Pos < 10'd100)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd480) && (X_Pos < 10'd485) && (Y_Pos > 10'd96) && (Y_Pos < 10'd100)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd96) && (Y_Pos < 10'd100)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd96) && (Y_Pos < 10'd100)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd97) && (Y_Pos < 10'd101)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd97) && (Y_Pos < 10'd101)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd154) && (X_Pos < 10'd159) && (Y_Pos > 10'd97) && (Y_Pos < 10'd101)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd97) && (Y_Pos < 10'd101)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd97) && (Y_Pos < 10'd101)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd280) && (X_Pos < 10'd285) && (Y_Pos > 10'd97) && (Y_Pos < 10'd101)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd97) && (Y_Pos < 10'd101)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd97) && (Y_Pos < 10'd101)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd354) && (X_Pos < 10'd359) && (Y_Pos > 10'd97) && (Y_Pos < 10'd101)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd97) && (Y_Pos < 10'd101)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd97) && (Y_Pos < 10'd101)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd480) && (X_Pos < 10'd485) && (Y_Pos > 10'd97) && (Y_Pos < 10'd101)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd97) && (Y_Pos < 10'd101)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd97) && (Y_Pos < 10'd101)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd98) && (Y_Pos < 10'd102)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd98) && (Y_Pos < 10'd102)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd154) && (X_Pos < 10'd159) && (Y_Pos > 10'd98) && (Y_Pos < 10'd102)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd98) && (Y_Pos < 10'd102)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd98) && (Y_Pos < 10'd102)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd280) && (X_Pos < 10'd285) && (Y_Pos > 10'd98) && (Y_Pos < 10'd102)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd98) && (Y_Pos < 10'd102)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd98) && (Y_Pos < 10'd102)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd354) && (X_Pos < 10'd359) && (Y_Pos > 10'd98) && (Y_Pos < 10'd102)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd98) && (Y_Pos < 10'd102)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd98) && (Y_Pos < 10'd102)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd480) && (X_Pos < 10'd485) && (Y_Pos > 10'd98) && (Y_Pos < 10'd102)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd98) && (Y_Pos < 10'd102)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd98) && (Y_Pos < 10'd102)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd99) && (Y_Pos < 10'd103)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd99) && (Y_Pos < 10'd103)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd154) && (X_Pos < 10'd159) && (Y_Pos > 10'd99) && (Y_Pos < 10'd103)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd99) && (Y_Pos < 10'd103)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd99) && (Y_Pos < 10'd103)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd280) && (X_Pos < 10'd285) && (Y_Pos > 10'd99) && (Y_Pos < 10'd103)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd99) && (Y_Pos < 10'd103)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd99) && (Y_Pos < 10'd103)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd354) && (X_Pos < 10'd359) && (Y_Pos > 10'd99) && (Y_Pos < 10'd103)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd99) && (Y_Pos < 10'd103)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd99) && (Y_Pos < 10'd103)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd480) && (X_Pos < 10'd485) && (Y_Pos > 10'd99) && (Y_Pos < 10'd103)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd99) && (Y_Pos < 10'd103)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd99) && (Y_Pos < 10'd103)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd100) && (Y_Pos < 10'd104)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd100) && (Y_Pos < 10'd104)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd154) && (X_Pos < 10'd159) && (Y_Pos > 10'd100) && (Y_Pos < 10'd104)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd194) && (X_Pos < 10'd199) && (Y_Pos > 10'd100) && (Y_Pos < 10'd104)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd100) && (Y_Pos < 10'd104)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd280) && (X_Pos < 10'd285) && (Y_Pos > 10'd100) && (Y_Pos < 10'd104)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd100) && (Y_Pos < 10'd104)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd100) && (Y_Pos < 10'd104)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd354) && (X_Pos < 10'd359) && (Y_Pos > 10'd100) && (Y_Pos < 10'd104)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd100) && (Y_Pos < 10'd104)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd440) && (X_Pos < 10'd445) && (Y_Pos > 10'd100) && (Y_Pos < 10'd104)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd480) && (X_Pos < 10'd485) && (Y_Pos > 10'd100) && (Y_Pos < 10'd104)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd100) && (Y_Pos < 10'd104)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd100) && (Y_Pos < 10'd104)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd101) && (Y_Pos < 10'd105)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd101) && (Y_Pos < 10'd105)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd155) && (X_Pos < 10'd160) && (Y_Pos > 10'd101) && (Y_Pos < 10'd105)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd193) && (X_Pos < 10'd198) && (Y_Pos > 10'd101) && (Y_Pos < 10'd105)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd227) && (X_Pos < 10'd232) && (Y_Pos > 10'd101) && (Y_Pos < 10'd105)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd279) && (X_Pos < 10'd284) && (Y_Pos > 10'd101) && (Y_Pos < 10'd105)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd312) && (X_Pos < 10'd318) && (Y_Pos > 10'd101) && (Y_Pos < 10'd105)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd321) && (X_Pos < 10'd327) && (Y_Pos > 10'd101) && (Y_Pos < 10'd105)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd355) && (X_Pos < 10'd360) && (Y_Pos > 10'd101) && (Y_Pos < 10'd105)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd407) && (X_Pos < 10'd412) && (Y_Pos > 10'd101) && (Y_Pos < 10'd105)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd441) && (X_Pos < 10'd446) && (Y_Pos > 10'd101) && (Y_Pos < 10'd105)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd479) && (X_Pos < 10'd484) && (Y_Pos > 10'd101) && (Y_Pos < 10'd105)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd101) && (Y_Pos < 10'd105)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd101) && (Y_Pos < 10'd105)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd102) && (Y_Pos < 10'd106)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd102) && (Y_Pos < 10'd106)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd156) && (X_Pos < 10'd197) && (Y_Pos > 10'd102) && (Y_Pos < 10'd106)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd227) && (X_Pos < 10'd283) && (Y_Pos > 10'd102) && (Y_Pos < 10'd106)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd313) && (X_Pos < 10'd326) && (Y_Pos > 10'd102) && (Y_Pos < 10'd106)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd356) && (X_Pos < 10'd412) && (Y_Pos > 10'd102) && (Y_Pos < 10'd106)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd442) && (X_Pos < 10'd483) && (Y_Pos > 10'd102) && (Y_Pos < 10'd106)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd102) && (Y_Pos < 10'd106)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd102) && (Y_Pos < 10'd106)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd103) && (Y_Pos < 10'd107)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd103) && (Y_Pos < 10'd107)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd157) && (X_Pos < 10'd196) && (Y_Pos > 10'd103) && (Y_Pos < 10'd107)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd229) && (X_Pos < 10'd282) && (Y_Pos > 10'd103) && (Y_Pos < 10'd107)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd315) && (X_Pos < 10'd324) && (Y_Pos > 10'd103) && (Y_Pos < 10'd107)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd357) && (X_Pos < 10'd410) && (Y_Pos > 10'd103) && (Y_Pos < 10'd107)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd443) && (X_Pos < 10'd482) && (Y_Pos > 10'd103) && (Y_Pos < 10'd107)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd103) && (Y_Pos < 10'd107)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd103) && (Y_Pos < 10'd107)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd104) && (Y_Pos < 10'd108)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd104) && (Y_Pos < 10'd108)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd104) && (Y_Pos < 10'd108)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd104) && (Y_Pos < 10'd108)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd105) && (Y_Pos < 10'd109)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd105) && (Y_Pos < 10'd109)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd105) && (Y_Pos < 10'd109)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd105) && (Y_Pos < 10'd109)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd106) && (Y_Pos < 10'd110)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd106) && (Y_Pos < 10'd110)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd106) && (Y_Pos < 10'd110)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd106) && (Y_Pos < 10'd110)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd107) && (Y_Pos < 10'd111)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd107) && (Y_Pos < 10'd111)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd107) && (Y_Pos < 10'd111)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd107) && (Y_Pos < 10'd111)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd108) && (Y_Pos < 10'd112)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd108) && (Y_Pos < 10'd112)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd108) && (Y_Pos < 10'd112)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd108) && (Y_Pos < 10'd112)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd109) && (Y_Pos < 10'd113)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd109) && (Y_Pos < 10'd113)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd109) && (Y_Pos < 10'd113)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd109) && (Y_Pos < 10'd113)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd110) && (Y_Pos < 10'd114)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd110) && (Y_Pos < 10'd114)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd110) && (Y_Pos < 10'd114)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd110) && (Y_Pos < 10'd114)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd111) && (Y_Pos < 10'd115)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd111) && (Y_Pos < 10'd115)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd111) && (Y_Pos < 10'd115)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd111) && (Y_Pos < 10'd115)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd112) && (Y_Pos < 10'd116)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd112) && (Y_Pos < 10'd116)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd112) && (Y_Pos < 10'd116)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd112) && (Y_Pos < 10'd116)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd113) && (Y_Pos < 10'd117)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd113) && (Y_Pos < 10'd117)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd113) && (Y_Pos < 10'd117)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd113) && (Y_Pos < 10'd117)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd114) && (Y_Pos < 10'd118)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd114) && (Y_Pos < 10'd118)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd114) && (Y_Pos < 10'd118)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd114) && (Y_Pos < 10'd118)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd115) && (Y_Pos < 10'd119)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd115) && (Y_Pos < 10'd119)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd115) && (Y_Pos < 10'd119)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd115) && (Y_Pos < 10'd119)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd116) && (Y_Pos < 10'd120)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd116) && (Y_Pos < 10'd120)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd116) && (Y_Pos < 10'd120)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd116) && (Y_Pos < 10'd120)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd117) && (Y_Pos < 10'd121)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd117) && (Y_Pos < 10'd121)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd117) && (Y_Pos < 10'd121)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd117) && (Y_Pos < 10'd121)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd118) && (Y_Pos < 10'd122)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd118) && (Y_Pos < 10'd122)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd118) && (Y_Pos < 10'd122)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd118) && (Y_Pos < 10'd122)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd119) && (Y_Pos < 10'd123)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd119) && (Y_Pos < 10'd123)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd119) && (Y_Pos < 10'd123)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd119) && (Y_Pos < 10'd123)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd120) && (Y_Pos < 10'd124)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd120) && (Y_Pos < 10'd124)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd120) && (Y_Pos < 10'd124)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd120) && (Y_Pos < 10'd124)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd121) && (Y_Pos < 10'd125)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd121) && (Y_Pos < 10'd125)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd121) && (Y_Pos < 10'd125)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd121) && (Y_Pos < 10'd125)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd122) && (Y_Pos < 10'd126)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd122) && (Y_Pos < 10'd126)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd122) && (Y_Pos < 10'd126)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd122) && (Y_Pos < 10'd126)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd123) && (Y_Pos < 10'd127)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd123) && (Y_Pos < 10'd127)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd123) && (Y_Pos < 10'd127)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd123) && (Y_Pos < 10'd127)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd124) && (Y_Pos < 10'd128)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd124) && (Y_Pos < 10'd128)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd124) && (Y_Pos < 10'd128)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd124) && (Y_Pos < 10'd128)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd125) && (Y_Pos < 10'd129)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd125) && (Y_Pos < 10'd129)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd125) && (Y_Pos < 10'd129)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd125) && (Y_Pos < 10'd129)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd126) && (Y_Pos < 10'd130)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd126) && (Y_Pos < 10'd130)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd126) && (Y_Pos < 10'd130)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd126) && (Y_Pos < 10'd130)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd127) && (Y_Pos < 10'd131)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd127) && (Y_Pos < 10'd131)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd127) && (Y_Pos < 10'd131)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd127) && (Y_Pos < 10'd131)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd128) && (Y_Pos < 10'd132)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd128) && (Y_Pos < 10'd132)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd128) && (Y_Pos < 10'd132)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd128) && (Y_Pos < 10'd132)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd129) && (Y_Pos < 10'd133)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd129) && (Y_Pos < 10'd133)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd129) && (Y_Pos < 10'd133)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd129) && (Y_Pos < 10'd133)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd130) && (Y_Pos < 10'd134)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd130) && (Y_Pos < 10'd134)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd157) && (X_Pos < 10'd196) && (Y_Pos > 10'd130) && (Y_Pos < 10'd134)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd229) && (X_Pos < 10'd239) && (Y_Pos > 10'd130) && (Y_Pos < 10'd134)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd272) && (X_Pos < 10'd367) && (Y_Pos > 10'd130) && (Y_Pos < 10'd134)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd400) && (X_Pos < 10'd410) && (Y_Pos > 10'd130) && (Y_Pos < 10'd134)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd443) && (X_Pos < 10'd482) && (Y_Pos > 10'd130) && (Y_Pos < 10'd134)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd130) && (Y_Pos < 10'd134)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd130) && (Y_Pos < 10'd134)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd131) && (Y_Pos < 10'd135)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd131) && (Y_Pos < 10'd135)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd156) && (X_Pos < 10'd197) && (Y_Pos > 10'd131) && (Y_Pos < 10'd135)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd227) && (X_Pos < 10'd240) && (Y_Pos > 10'd131) && (Y_Pos < 10'd135)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd270) && (X_Pos < 10'd369) && (Y_Pos > 10'd131) && (Y_Pos < 10'd135)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd399) && (X_Pos < 10'd412) && (Y_Pos > 10'd131) && (Y_Pos < 10'd135)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd442) && (X_Pos < 10'd483) && (Y_Pos > 10'd131) && (Y_Pos < 10'd135)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd131) && (Y_Pos < 10'd135)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd131) && (Y_Pos < 10'd135)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd132) && (Y_Pos < 10'd136)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd132) && (Y_Pos < 10'd136)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd155) && (X_Pos < 10'd160) && (Y_Pos > 10'd132) && (Y_Pos < 10'd136)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd193) && (X_Pos < 10'd198) && (Y_Pos > 10'd132) && (Y_Pos < 10'd136)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd227) && (X_Pos < 10'd232) && (Y_Pos > 10'd132) && (Y_Pos < 10'd136)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd236) && (X_Pos < 10'd241) && (Y_Pos > 10'd132) && (Y_Pos < 10'd136)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd270) && (X_Pos < 10'd275) && (Y_Pos > 10'd132) && (Y_Pos < 10'd136)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd364) && (X_Pos < 10'd369) && (Y_Pos > 10'd132) && (Y_Pos < 10'd136)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd398) && (X_Pos < 10'd403) && (Y_Pos > 10'd132) && (Y_Pos < 10'd136)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd407) && (X_Pos < 10'd412) && (Y_Pos > 10'd132) && (Y_Pos < 10'd136)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd441) && (X_Pos < 10'd446) && (Y_Pos > 10'd132) && (Y_Pos < 10'd136)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd479) && (X_Pos < 10'd484) && (Y_Pos > 10'd132) && (Y_Pos < 10'd136)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd132) && (Y_Pos < 10'd136)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd132) && (Y_Pos < 10'd136)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd133) && (Y_Pos < 10'd137)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd133) && (Y_Pos < 10'd137)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd154) && (X_Pos < 10'd159) && (Y_Pos > 10'd133) && (Y_Pos < 10'd137)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd194) && (X_Pos < 10'd200) && (Y_Pos > 10'd133) && (Y_Pos < 10'd137)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd133) && (Y_Pos < 10'd137)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd237) && (X_Pos < 10'd242) && (Y_Pos > 10'd133) && (Y_Pos < 10'd137)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd133) && (Y_Pos < 10'd137)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd133) && (Y_Pos < 10'd137)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd397) && (X_Pos < 10'd402) && (Y_Pos > 10'd133) && (Y_Pos < 10'd137)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd133) && (Y_Pos < 10'd137)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd445) && (Y_Pos > 10'd133) && (Y_Pos < 10'd137)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd480) && (X_Pos < 10'd485) && (Y_Pos > 10'd133) && (Y_Pos < 10'd137)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd133) && (Y_Pos < 10'd137)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd133) && (Y_Pos < 10'd137)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd134) && (Y_Pos < 10'd138)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd134) && (Y_Pos < 10'd138)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd154) && (X_Pos < 10'd159) && (Y_Pos > 10'd134) && (Y_Pos < 10'd138)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd134) && (Y_Pos < 10'd138)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd134) && (Y_Pos < 10'd138)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd134) && (Y_Pos < 10'd138)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd134) && (Y_Pos < 10'd138)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd134) && (Y_Pos < 10'd138)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd134) && (Y_Pos < 10'd138)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd134) && (Y_Pos < 10'd138)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd134) && (Y_Pos < 10'd138)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd480) && (X_Pos < 10'd485) && (Y_Pos > 10'd134) && (Y_Pos < 10'd138)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd134) && (Y_Pos < 10'd138)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd134) && (Y_Pos < 10'd138)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd135) && (Y_Pos < 10'd139)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd135) && (Y_Pos < 10'd139)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd154) && (X_Pos < 10'd159) && (Y_Pos > 10'd135) && (Y_Pos < 10'd139)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd135) && (Y_Pos < 10'd139)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd135) && (Y_Pos < 10'd139)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd135) && (Y_Pos < 10'd139)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd135) && (Y_Pos < 10'd139)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd135) && (Y_Pos < 10'd139)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd135) && (Y_Pos < 10'd139)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd135) && (Y_Pos < 10'd139)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd135) && (Y_Pos < 10'd139)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd480) && (X_Pos < 10'd485) && (Y_Pos > 10'd135) && (Y_Pos < 10'd139)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd135) && (Y_Pos < 10'd139)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd135) && (Y_Pos < 10'd139)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd136) && (Y_Pos < 10'd140)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd136) && (Y_Pos < 10'd140)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd154) && (X_Pos < 10'd159) && (Y_Pos > 10'd136) && (Y_Pos < 10'd140)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd136) && (Y_Pos < 10'd140)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd136) && (Y_Pos < 10'd140)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd136) && (Y_Pos < 10'd140)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd136) && (Y_Pos < 10'd140)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd136) && (Y_Pos < 10'd140)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd136) && (Y_Pos < 10'd140)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd136) && (Y_Pos < 10'd140)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd136) && (Y_Pos < 10'd140)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd480) && (X_Pos < 10'd485) && (Y_Pos > 10'd136) && (Y_Pos < 10'd140)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd136) && (Y_Pos < 10'd140)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd136) && (Y_Pos < 10'd140)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd137) && (Y_Pos < 10'd141)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd137) && (Y_Pos < 10'd141)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd154) && (X_Pos < 10'd159) && (Y_Pos > 10'd137) && (Y_Pos < 10'd141)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd137) && (Y_Pos < 10'd141)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd137) && (Y_Pos < 10'd141)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd137) && (Y_Pos < 10'd141)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd137) && (Y_Pos < 10'd141)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd137) && (Y_Pos < 10'd141)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd137) && (Y_Pos < 10'd141)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd137) && (Y_Pos < 10'd141)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd137) && (Y_Pos < 10'd141)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd480) && (X_Pos < 10'd485) && (Y_Pos > 10'd137) && (Y_Pos < 10'd141)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd137) && (Y_Pos < 10'd141)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd137) && (Y_Pos < 10'd141)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd138) && (Y_Pos < 10'd142)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd138) && (Y_Pos < 10'd142)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd154) && (X_Pos < 10'd159) && (Y_Pos > 10'd138) && (Y_Pos < 10'd142)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd138) && (Y_Pos < 10'd142)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd138) && (Y_Pos < 10'd142)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd138) && (Y_Pos < 10'd142)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd138) && (Y_Pos < 10'd142)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd138) && (Y_Pos < 10'd142)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd138) && (Y_Pos < 10'd142)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd138) && (Y_Pos < 10'd142)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd138) && (Y_Pos < 10'd142)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd480) && (X_Pos < 10'd485) && (Y_Pos > 10'd138) && (Y_Pos < 10'd142)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd138) && (Y_Pos < 10'd142)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd138) && (Y_Pos < 10'd142)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd139) && (Y_Pos < 10'd143)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd139) && (Y_Pos < 10'd143)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd154) && (X_Pos < 10'd160) && (Y_Pos > 10'd139) && (Y_Pos < 10'd143)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd194) && (X_Pos < 10'd199) && (Y_Pos > 10'd139) && (Y_Pos < 10'd143)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd139) && (Y_Pos < 10'd143)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd139) && (Y_Pos < 10'd143)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd269) && (X_Pos < 10'd274) && (Y_Pos > 10'd139) && (Y_Pos < 10'd143)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd365) && (X_Pos < 10'd370) && (Y_Pos > 10'd139) && (Y_Pos < 10'd143)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd139) && (Y_Pos < 10'd143)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd139) && (Y_Pos < 10'd143)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd440) && (X_Pos < 10'd445) && (Y_Pos > 10'd139) && (Y_Pos < 10'd143)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd479) && (X_Pos < 10'd485) && (Y_Pos > 10'd139) && (Y_Pos < 10'd143)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd139) && (Y_Pos < 10'd143)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd139) && (Y_Pos < 10'd143)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd140) && (Y_Pos < 10'd144)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd140) && (Y_Pos < 10'd144)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd155) && (X_Pos < 10'd160) && (Y_Pos > 10'd140) && (Y_Pos < 10'd144)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd193) && (X_Pos < 10'd198) && (Y_Pos > 10'd140) && (Y_Pos < 10'd144)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd140) && (Y_Pos < 10'd144)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd140) && (Y_Pos < 10'd144)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd270) && (X_Pos < 10'd275) && (Y_Pos > 10'd140) && (Y_Pos < 10'd144)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd364) && (X_Pos < 10'd369) && (Y_Pos > 10'd140) && (Y_Pos < 10'd144)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd140) && (Y_Pos < 10'd144)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd140) && (Y_Pos < 10'd144)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd441) && (X_Pos < 10'd446) && (Y_Pos > 10'd140) && (Y_Pos < 10'd144)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd479) && (X_Pos < 10'd484) && (Y_Pos > 10'd140) && (Y_Pos < 10'd144)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd140) && (Y_Pos < 10'd144)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd140) && (Y_Pos < 10'd144)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd141) && (Y_Pos < 10'd145)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd141) && (Y_Pos < 10'd145)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd157) && (X_Pos < 10'd196) && (Y_Pos > 10'd141) && (Y_Pos < 10'd145)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd141) && (Y_Pos < 10'd145)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd141) && (Y_Pos < 10'd145)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd271) && (X_Pos < 10'd312) && (Y_Pos > 10'd141) && (Y_Pos < 10'd145)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd327) && (X_Pos < 10'd368) && (Y_Pos > 10'd141) && (Y_Pos < 10'd145)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd141) && (Y_Pos < 10'd145)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd141) && (Y_Pos < 10'd145)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd443) && (X_Pos < 10'd482) && (Y_Pos > 10'd141) && (Y_Pos < 10'd145)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd141) && (Y_Pos < 10'd145)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd141) && (Y_Pos < 10'd145)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd142) && (Y_Pos < 10'd146)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd142) && (Y_Pos < 10'd146)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd158) && (X_Pos < 10'd196) && (Y_Pos > 10'd142) && (Y_Pos < 10'd146)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd142) && (Y_Pos < 10'd146)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd142) && (Y_Pos < 10'd146)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd272) && (X_Pos < 10'd313) && (Y_Pos > 10'd142) && (Y_Pos < 10'd146)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd326) && (X_Pos < 10'd367) && (Y_Pos > 10'd142) && (Y_Pos < 10'd146)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd142) && (Y_Pos < 10'd146)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd142) && (Y_Pos < 10'd146)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd443) && (X_Pos < 10'd481) && (Y_Pos > 10'd142) && (Y_Pos < 10'd146)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd142) && (Y_Pos < 10'd146)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd142) && (Y_Pos < 10'd146)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd143) && (Y_Pos < 10'd147)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd143) && (Y_Pos < 10'd147)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd143) && (Y_Pos < 10'd147)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd143) && (Y_Pos < 10'd147)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd309) && (X_Pos < 10'd314) && (Y_Pos > 10'd143) && (Y_Pos < 10'd147)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd325) && (X_Pos < 10'd330) && (Y_Pos > 10'd143) && (Y_Pos < 10'd147)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd143) && (Y_Pos < 10'd147)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd143) && (Y_Pos < 10'd147)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd143) && (Y_Pos < 10'd147)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd143) && (Y_Pos < 10'd147)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd144) && (Y_Pos < 10'd148)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd144) && (Y_Pos < 10'd148)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd144) && (Y_Pos < 10'd148)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd144) && (Y_Pos < 10'd148)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd310) && (X_Pos < 10'd315) && (Y_Pos > 10'd144) && (Y_Pos < 10'd148)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd324) && (X_Pos < 10'd329) && (Y_Pos > 10'd144) && (Y_Pos < 10'd148)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd144) && (Y_Pos < 10'd148)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd144) && (Y_Pos < 10'd148)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd144) && (Y_Pos < 10'd148)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd144) && (Y_Pos < 10'd148)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd145) && (Y_Pos < 10'd149)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd145) && (Y_Pos < 10'd149)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd145) && (Y_Pos < 10'd149)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd145) && (Y_Pos < 10'd149)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd145) && (Y_Pos < 10'd149)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd145) && (Y_Pos < 10'd149)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd145) && (Y_Pos < 10'd149)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd145) && (Y_Pos < 10'd149)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd145) && (Y_Pos < 10'd149)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd145) && (Y_Pos < 10'd149)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd146) && (Y_Pos < 10'd150)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd146) && (Y_Pos < 10'd150)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd146) && (Y_Pos < 10'd150)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd146) && (Y_Pos < 10'd150)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd146) && (Y_Pos < 10'd150)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd146) && (Y_Pos < 10'd150)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd146) && (Y_Pos < 10'd150)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd146) && (Y_Pos < 10'd150)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd146) && (Y_Pos < 10'd150)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd146) && (Y_Pos < 10'd150)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd147) && (Y_Pos < 10'd151)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd147) && (Y_Pos < 10'd151)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd147) && (Y_Pos < 10'd151)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd147) && (Y_Pos < 10'd151)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd147) && (Y_Pos < 10'd151)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd147) && (Y_Pos < 10'd151)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd147) && (Y_Pos < 10'd151)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd147) && (Y_Pos < 10'd151)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd147) && (Y_Pos < 10'd151)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd147) && (Y_Pos < 10'd151)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd148) && (Y_Pos < 10'd152)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd148) && (Y_Pos < 10'd152)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd148) && (Y_Pos < 10'd152)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd148) && (Y_Pos < 10'd152)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd148) && (Y_Pos < 10'd152)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd148) && (Y_Pos < 10'd152)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd148) && (Y_Pos < 10'd152)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd148) && (Y_Pos < 10'd152)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd148) && (Y_Pos < 10'd152)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd148) && (Y_Pos < 10'd152)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd149) && (Y_Pos < 10'd153)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd149) && (Y_Pos < 10'd153)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd149) && (Y_Pos < 10'd153)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd149) && (Y_Pos < 10'd153)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd149) && (Y_Pos < 10'd153)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd149) && (Y_Pos < 10'd153)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd149) && (Y_Pos < 10'd153)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd149) && (Y_Pos < 10'd153)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd149) && (Y_Pos < 10'd153)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd149) && (Y_Pos < 10'd153)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd150) && (Y_Pos < 10'd154)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd150) && (Y_Pos < 10'd154)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd150) && (Y_Pos < 10'd154)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd150) && (Y_Pos < 10'd154)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd150) && (Y_Pos < 10'd154)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd150) && (Y_Pos < 10'd154)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd150) && (Y_Pos < 10'd154)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd150) && (Y_Pos < 10'd154)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd150) && (Y_Pos < 10'd154)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd150) && (Y_Pos < 10'd154)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd151) && (Y_Pos < 10'd155)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd151) && (Y_Pos < 10'd155)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd151) && (Y_Pos < 10'd155)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd151) && (Y_Pos < 10'd155)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd151) && (Y_Pos < 10'd155)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd151) && (Y_Pos < 10'd155)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd151) && (Y_Pos < 10'd155)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd151) && (Y_Pos < 10'd155)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd151) && (Y_Pos < 10'd155)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd151) && (Y_Pos < 10'd155)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd152) && (Y_Pos < 10'd156)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd152) && (Y_Pos < 10'd156)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd152) && (Y_Pos < 10'd156)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd152) && (Y_Pos < 10'd156)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd152) && (Y_Pos < 10'd156)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd152) && (Y_Pos < 10'd156)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd152) && (Y_Pos < 10'd156)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd152) && (Y_Pos < 10'd156)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd152) && (Y_Pos < 10'd156)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd152) && (Y_Pos < 10'd156)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd153) && (Y_Pos < 10'd157)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd153) && (Y_Pos < 10'd157)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd153) && (Y_Pos < 10'd157)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd153) && (Y_Pos < 10'd157)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd153) && (Y_Pos < 10'd157)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd153) && (Y_Pos < 10'd157)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd153) && (Y_Pos < 10'd157)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd153) && (Y_Pos < 10'd157)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd153) && (Y_Pos < 10'd157)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd153) && (Y_Pos < 10'd157)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd154) && (Y_Pos < 10'd158)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd154) && (Y_Pos < 10'd158)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd154) && (Y_Pos < 10'd158)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd154) && (Y_Pos < 10'd158)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd154) && (Y_Pos < 10'd158)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd154) && (Y_Pos < 10'd158)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd154) && (Y_Pos < 10'd158)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd154) && (Y_Pos < 10'd158)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd154) && (Y_Pos < 10'd158)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd154) && (Y_Pos < 10'd158)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd155) && (Y_Pos < 10'd159)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd155) && (Y_Pos < 10'd159)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd155) && (Y_Pos < 10'd159)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd155) && (Y_Pos < 10'd159)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd155) && (Y_Pos < 10'd159)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd155) && (Y_Pos < 10'd159)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd155) && (Y_Pos < 10'd159)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd155) && (Y_Pos < 10'd159)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd155) && (Y_Pos < 10'd159)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd155) && (Y_Pos < 10'd159)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd156) && (Y_Pos < 10'd160)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd156) && (Y_Pos < 10'd160)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd156) && (Y_Pos < 10'd160)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd156) && (Y_Pos < 10'd160)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd156) && (Y_Pos < 10'd160)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd156) && (Y_Pos < 10'd160)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd156) && (Y_Pos < 10'd160)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd156) && (Y_Pos < 10'd160)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd156) && (Y_Pos < 10'd160)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd156) && (Y_Pos < 10'd160)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd157) && (Y_Pos < 10'd161)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd157) && (Y_Pos < 10'd161)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd157) && (Y_Pos < 10'd161)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd157) && (Y_Pos < 10'd161)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd157) && (Y_Pos < 10'd161)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd157) && (Y_Pos < 10'd161)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd157) && (Y_Pos < 10'd161)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd157) && (Y_Pos < 10'd161)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd157) && (Y_Pos < 10'd161)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd157) && (Y_Pos < 10'd161)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd158) && (Y_Pos < 10'd162)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd158) && (Y_Pos < 10'd162)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd158) && (Y_Pos < 10'd162)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd158) && (Y_Pos < 10'd162)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd158) && (Y_Pos < 10'd162)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd158) && (Y_Pos < 10'd162)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd158) && (Y_Pos < 10'd162)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd158) && (Y_Pos < 10'd162)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd158) && (Y_Pos < 10'd162)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd158) && (Y_Pos < 10'd162)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd159) && (Y_Pos < 10'd163)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd159) && (Y_Pos < 10'd163)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd159) && (Y_Pos < 10'd163)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd159) && (Y_Pos < 10'd163)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd159) && (Y_Pos < 10'd163)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd159) && (Y_Pos < 10'd163)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd159) && (Y_Pos < 10'd163)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd159) && (Y_Pos < 10'd163)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd159) && (Y_Pos < 10'd163)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd159) && (Y_Pos < 10'd163)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd160) && (Y_Pos < 10'd164)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd160) && (Y_Pos < 10'd164)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd160) && (Y_Pos < 10'd164)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd160) && (Y_Pos < 10'd164)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd160) && (Y_Pos < 10'd164)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd160) && (Y_Pos < 10'd164)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd160) && (Y_Pos < 10'd164)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd160) && (Y_Pos < 10'd164)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd160) && (Y_Pos < 10'd164)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd160) && (Y_Pos < 10'd164)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd161) && (Y_Pos < 10'd165)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd161) && (Y_Pos < 10'd165)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd161) && (Y_Pos < 10'd165)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd161) && (Y_Pos < 10'd165)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd161) && (Y_Pos < 10'd165)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd161) && (Y_Pos < 10'd165)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd161) && (Y_Pos < 10'd165)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd161) && (Y_Pos < 10'd165)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd161) && (Y_Pos < 10'd165)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd161) && (Y_Pos < 10'd165)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd162) && (Y_Pos < 10'd166)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd162) && (Y_Pos < 10'd166)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd162) && (Y_Pos < 10'd166)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd162) && (Y_Pos < 10'd166)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd162) && (Y_Pos < 10'd166)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd162) && (Y_Pos < 10'd166)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd162) && (Y_Pos < 10'd166)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd162) && (Y_Pos < 10'd166)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd162) && (Y_Pos < 10'd166)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd162) && (Y_Pos < 10'd166)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd163) && (Y_Pos < 10'd167)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd163) && (Y_Pos < 10'd167)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd163) && (Y_Pos < 10'd167)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd163) && (Y_Pos < 10'd167)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd163) && (Y_Pos < 10'd167)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd163) && (Y_Pos < 10'd167)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd163) && (Y_Pos < 10'd167)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd163) && (Y_Pos < 10'd167)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd163) && (Y_Pos < 10'd167)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd163) && (Y_Pos < 10'd167)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd164) && (Y_Pos < 10'd168)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd164) && (Y_Pos < 10'd168)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd164) && (Y_Pos < 10'd168)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd164) && (Y_Pos < 10'd168)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd164) && (Y_Pos < 10'd168)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd164) && (Y_Pos < 10'd168)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd164) && (Y_Pos < 10'd168)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd164) && (Y_Pos < 10'd168)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd164) && (Y_Pos < 10'd168)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd164) && (Y_Pos < 10'd168)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd165) && (Y_Pos < 10'd169)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd165) && (Y_Pos < 10'd169)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd165) && (Y_Pos < 10'd169)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd237) && (X_Pos < 10'd243) && (Y_Pos > 10'd165) && (Y_Pos < 10'd169)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd165) && (Y_Pos < 10'd169)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd165) && (Y_Pos < 10'd169)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd402) && (Y_Pos > 10'd165) && (Y_Pos < 10'd169)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd165) && (Y_Pos < 10'd169)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd165) && (Y_Pos < 10'd169)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd165) && (Y_Pos < 10'd169)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd166) && (Y_Pos < 10'd170)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd166) && (Y_Pos < 10'd170)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd166) && (Y_Pos < 10'd170)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd166) && (Y_Pos < 10'd170)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd166) && (Y_Pos < 10'd170)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd166) && (Y_Pos < 10'd170)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd166) && (Y_Pos < 10'd170)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd166) && (Y_Pos < 10'd170)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd166) && (Y_Pos < 10'd170)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd166) && (Y_Pos < 10'd170)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd167) && (Y_Pos < 10'd171)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd125) && (X_Pos < 10'd130) && (Y_Pos > 10'd167) && (Y_Pos < 10'd171)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd167) && (Y_Pos < 10'd171)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd239) && (X_Pos < 10'd244) && (Y_Pos > 10'd167) && (Y_Pos < 10'd171)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd167) && (Y_Pos < 10'd171)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd167) && (Y_Pos < 10'd171)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd395) && (X_Pos < 10'd400) && (Y_Pos > 10'd167) && (Y_Pos < 10'd171)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd167) && (Y_Pos < 10'd171)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd509) && (X_Pos < 10'd514) && (Y_Pos > 10'd167) && (Y_Pos < 10'd171)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd167) && (Y_Pos < 10'd171)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd168) && (Y_Pos < 10'd172)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd125) && (X_Pos < 10'd195) && (Y_Pos > 10'd168) && (Y_Pos < 10'd172)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd168) && (Y_Pos < 10'd172)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd240) && (X_Pos < 10'd281) && (Y_Pos > 10'd168) && (Y_Pos < 10'd172)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd168) && (Y_Pos < 10'd172)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd168) && (Y_Pos < 10'd172)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd358) && (X_Pos < 10'd399) && (Y_Pos > 10'd168) && (Y_Pos < 10'd172)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd168) && (Y_Pos < 10'd172)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd444) && (X_Pos < 10'd514) && (Y_Pos > 10'd168) && (Y_Pos < 10'd172)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd168) && (Y_Pos < 10'd172)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd120) && (X_Pos < 10'd125) && (Y_Pos > 10'd169) && (Y_Pos < 10'd173)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd127) && (X_Pos < 10'd196) && (Y_Pos > 10'd169) && (Y_Pos < 10'd173)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd169) && (Y_Pos < 10'd173)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd241) && (X_Pos < 10'd282) && (Y_Pos > 10'd169) && (Y_Pos < 10'd173)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd169) && (Y_Pos < 10'd173)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd169) && (Y_Pos < 10'd173)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd357) && (X_Pos < 10'd398) && (Y_Pos > 10'd169) && (Y_Pos < 10'd173)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd169) && (Y_Pos < 10'd173)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd443) && (X_Pos < 10'd512) && (Y_Pos > 10'd169) && (Y_Pos < 10'd173)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd514) && (X_Pos < 10'd519) && (Y_Pos > 10'd169) && (Y_Pos < 10'd173)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd120) && (X_Pos < 10'd125) && (Y_Pos > 10'd170) && (Y_Pos < 10'd174)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd193) && (X_Pos < 10'd198) && (Y_Pos > 10'd170) && (Y_Pos < 10'd174)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd170) && (Y_Pos < 10'd174)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd278) && (X_Pos < 10'd283) && (Y_Pos > 10'd170) && (Y_Pos < 10'd174)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd170) && (Y_Pos < 10'd174)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd170) && (Y_Pos < 10'd174)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd356) && (X_Pos < 10'd361) && (Y_Pos > 10'd170) && (Y_Pos < 10'd174)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd170) && (Y_Pos < 10'd174)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd441) && (X_Pos < 10'd446) && (Y_Pos > 10'd170) && (Y_Pos < 10'd174)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd514) && (X_Pos < 10'd519) && (Y_Pos > 10'd170) && (Y_Pos < 10'd174)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd120) && (X_Pos < 10'd125) && (Y_Pos > 10'd171) && (Y_Pos < 10'd175)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd193) && (X_Pos < 10'd198) && (Y_Pos > 10'd171) && (Y_Pos < 10'd175)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd171) && (Y_Pos < 10'd175)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd279) && (X_Pos < 10'd284) && (Y_Pos > 10'd171) && (Y_Pos < 10'd175)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd171) && (Y_Pos < 10'd175)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd171) && (Y_Pos < 10'd175)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd355) && (X_Pos < 10'd360) && (Y_Pos > 10'd171) && (Y_Pos < 10'd175)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd171) && (Y_Pos < 10'd175)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd441) && (X_Pos < 10'd446) && (Y_Pos > 10'd171) && (Y_Pos < 10'd175)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd514) && (X_Pos < 10'd519) && (Y_Pos > 10'd171) && (Y_Pos < 10'd175)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd122) && (X_Pos < 10'd128) && (Y_Pos > 10'd172) && (Y_Pos < 10'd176)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd172) && (Y_Pos < 10'd176)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd172) && (Y_Pos < 10'd176)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd280) && (X_Pos < 10'd285) && (Y_Pos > 10'd172) && (Y_Pos < 10'd176)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd172) && (Y_Pos < 10'd176)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd172) && (Y_Pos < 10'd176)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd354) && (X_Pos < 10'd359) && (Y_Pos > 10'd172) && (Y_Pos < 10'd176)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd172) && (Y_Pos < 10'd176)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd172) && (Y_Pos < 10'd176)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd517) && (Y_Pos > 10'd172) && (Y_Pos < 10'd176)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd122) && (X_Pos < 10'd192) && (Y_Pos > 10'd173) && (Y_Pos < 10'd177)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd173) && (Y_Pos < 10'd177)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd173) && (Y_Pos < 10'd177)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd280) && (X_Pos < 10'd285) && (Y_Pos > 10'd173) && (Y_Pos < 10'd177)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd173) && (Y_Pos < 10'd177)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd173) && (Y_Pos < 10'd177)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd354) && (X_Pos < 10'd359) && (Y_Pos > 10'd173) && (Y_Pos < 10'd177)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd173) && (Y_Pos < 10'd177)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd173) && (Y_Pos < 10'd177)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd447) && (X_Pos < 10'd517) && (Y_Pos > 10'd173) && (Y_Pos < 10'd177)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd125) && (X_Pos < 10'd193) && (Y_Pos > 10'd174) && (Y_Pos < 10'd178)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd174) && (Y_Pos < 10'd178)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd174) && (Y_Pos < 10'd178)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd280) && (X_Pos < 10'd285) && (Y_Pos > 10'd174) && (Y_Pos < 10'd178)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd174) && (Y_Pos < 10'd178)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd174) && (Y_Pos < 10'd178)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd354) && (X_Pos < 10'd359) && (Y_Pos > 10'd174) && (Y_Pos < 10'd178)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd174) && (Y_Pos < 10'd178)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd174) && (Y_Pos < 10'd178)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd446) && (X_Pos < 10'd514) && (Y_Pos > 10'd174) && (Y_Pos < 10'd178)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd175) && (Y_Pos < 10'd179)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd175) && (Y_Pos < 10'd179)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd175) && (Y_Pos < 10'd179)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd280) && (X_Pos < 10'd285) && (Y_Pos > 10'd175) && (Y_Pos < 10'd179)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd175) && (Y_Pos < 10'd179)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd175) && (Y_Pos < 10'd179)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd354) && (X_Pos < 10'd359) && (Y_Pos > 10'd175) && (Y_Pos < 10'd179)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd175) && (Y_Pos < 10'd179)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd175) && (Y_Pos < 10'd179)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd175) && (Y_Pos < 10'd179)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd176) && (Y_Pos < 10'd180)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd176) && (Y_Pos < 10'd180)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd176) && (Y_Pos < 10'd180)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd280) && (X_Pos < 10'd285) && (Y_Pos > 10'd176) && (Y_Pos < 10'd180)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd176) && (Y_Pos < 10'd180)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd176) && (Y_Pos < 10'd180)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd354) && (X_Pos < 10'd359) && (Y_Pos > 10'd176) && (Y_Pos < 10'd180)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd176) && (Y_Pos < 10'd180)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd176) && (Y_Pos < 10'd180)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd176) && (Y_Pos < 10'd180)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd177) && (Y_Pos < 10'd181)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd177) && (Y_Pos < 10'd181)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd177) && (Y_Pos < 10'd181)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd280) && (X_Pos < 10'd285) && (Y_Pos > 10'd177) && (Y_Pos < 10'd181)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd177) && (Y_Pos < 10'd181)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd177) && (Y_Pos < 10'd181)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd354) && (X_Pos < 10'd359) && (Y_Pos > 10'd177) && (Y_Pos < 10'd181)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd177) && (Y_Pos < 10'd181)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd177) && (Y_Pos < 10'd181)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd177) && (Y_Pos < 10'd181)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd178) && (Y_Pos < 10'd182)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd178) && (Y_Pos < 10'd182)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd178) && (Y_Pos < 10'd182)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd279) && (X_Pos < 10'd284) && (Y_Pos > 10'd178) && (Y_Pos < 10'd182)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd312) && (X_Pos < 10'd317) && (Y_Pos > 10'd178) && (Y_Pos < 10'd182)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd322) && (X_Pos < 10'd327) && (Y_Pos > 10'd178) && (Y_Pos < 10'd182)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd355) && (X_Pos < 10'd360) && (Y_Pos > 10'd178) && (Y_Pos < 10'd182)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd178) && (Y_Pos < 10'd182)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd178) && (Y_Pos < 10'd182)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd178) && (Y_Pos < 10'd182)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd179) && (Y_Pos < 10'd183)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd179) && (Y_Pos < 10'd183)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd179) && (Y_Pos < 10'd183)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd278) && (X_Pos < 10'd283) && (Y_Pos > 10'd179) && (Y_Pos < 10'd183)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd313) && (X_Pos < 10'd318) && (Y_Pos > 10'd179) && (Y_Pos < 10'd183)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd321) && (X_Pos < 10'd326) && (Y_Pos > 10'd179) && (Y_Pos < 10'd183)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd356) && (X_Pos < 10'd361) && (Y_Pos > 10'd179) && (Y_Pos < 10'd183)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd179) && (Y_Pos < 10'd183)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd179) && (Y_Pos < 10'd183)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd179) && (Y_Pos < 10'd183)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd180) && (Y_Pos < 10'd184)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd180) && (Y_Pos < 10'd184)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd180) && (Y_Pos < 10'd184)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd241) && (X_Pos < 10'd282) && (Y_Pos > 10'd180) && (Y_Pos < 10'd184)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd314) && (X_Pos < 10'd325) && (Y_Pos > 10'd180) && (Y_Pos < 10'd184)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd357) && (X_Pos < 10'd398) && (Y_Pos > 10'd180) && (Y_Pos < 10'd184)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd180) && (Y_Pos < 10'd184)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd180) && (Y_Pos < 10'd184)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd180) && (Y_Pos < 10'd184)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd181) && (Y_Pos < 10'd185)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd181) && (Y_Pos < 10'd185)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd181) && (Y_Pos < 10'd185)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd240) && (X_Pos < 10'd281) && (Y_Pos > 10'd181) && (Y_Pos < 10'd185)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd315) && (X_Pos < 10'd324) && (Y_Pos > 10'd181) && (Y_Pos < 10'd185)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd358) && (X_Pos < 10'd399) && (Y_Pos > 10'd181) && (Y_Pos < 10'd185)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd181) && (Y_Pos < 10'd185)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd181) && (Y_Pos < 10'd185)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd181) && (Y_Pos < 10'd185)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd182) && (Y_Pos < 10'd186)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd182) && (Y_Pos < 10'd186)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd182) && (Y_Pos < 10'd186)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd239) && (X_Pos < 10'd244) && (Y_Pos > 10'd182) && (Y_Pos < 10'd186)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd395) && (X_Pos < 10'd400) && (Y_Pos > 10'd182) && (Y_Pos < 10'd186)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd182) && (Y_Pos < 10'd186)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd182) && (Y_Pos < 10'd186)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd182) && (Y_Pos < 10'd186)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd183) && (Y_Pos < 10'd187)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd183) && (Y_Pos < 10'd187)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd183) && (Y_Pos < 10'd187)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd183) && (Y_Pos < 10'd187)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd183) && (Y_Pos < 10'd187)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd183) && (Y_Pos < 10'd187)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd183) && (Y_Pos < 10'd187)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd183) && (Y_Pos < 10'd187)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd184) && (Y_Pos < 10'd188)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd184) && (Y_Pos < 10'd188)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd184) && (Y_Pos < 10'd188)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd237) && (X_Pos < 10'd243) && (Y_Pos > 10'd184) && (Y_Pos < 10'd188)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd402) && (Y_Pos > 10'd184) && (Y_Pos < 10'd188)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd184) && (Y_Pos < 10'd188)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd184) && (Y_Pos < 10'd188)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd184) && (Y_Pos < 10'd188)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd185) && (Y_Pos < 10'd189)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd185) && (Y_Pos < 10'd189)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd185) && (Y_Pos < 10'd189)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd185) && (Y_Pos < 10'd189)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd185) && (Y_Pos < 10'd189)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd185) && (Y_Pos < 10'd189)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd185) && (Y_Pos < 10'd189)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd185) && (Y_Pos < 10'd189)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd186) && (Y_Pos < 10'd190)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd186) && (Y_Pos < 10'd190)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd186) && (Y_Pos < 10'd190)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd186) && (Y_Pos < 10'd190)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd186) && (Y_Pos < 10'd190)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd186) && (Y_Pos < 10'd190)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd186) && (Y_Pos < 10'd190)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd186) && (Y_Pos < 10'd190)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd187) && (Y_Pos < 10'd191)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd187) && (Y_Pos < 10'd191)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd187) && (Y_Pos < 10'd191)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd187) && (Y_Pos < 10'd191)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd187) && (Y_Pos < 10'd191)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd187) && (Y_Pos < 10'd191)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd187) && (Y_Pos < 10'd191)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd187) && (Y_Pos < 10'd191)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd188) && (Y_Pos < 10'd192)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd188) && (Y_Pos < 10'd192)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd188) && (Y_Pos < 10'd192)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd188) && (Y_Pos < 10'd192)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd188) && (Y_Pos < 10'd192)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd188) && (Y_Pos < 10'd192)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd188) && (Y_Pos < 10'd192)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd188) && (Y_Pos < 10'd192)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd189) && (Y_Pos < 10'd193)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd189) && (Y_Pos < 10'd193)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd189) && (Y_Pos < 10'd193)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd189) && (Y_Pos < 10'd193)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd189) && (Y_Pos < 10'd193)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd189) && (Y_Pos < 10'd193)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd189) && (Y_Pos < 10'd193)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd189) && (Y_Pos < 10'd193)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd190) && (Y_Pos < 10'd194)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd190) && (Y_Pos < 10'd194)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd190) && (Y_Pos < 10'd194)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd190) && (Y_Pos < 10'd194)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd190) && (Y_Pos < 10'd194)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd190) && (Y_Pos < 10'd194)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd190) && (Y_Pos < 10'd194)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd190) && (Y_Pos < 10'd194)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd191) && (Y_Pos < 10'd195)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd191) && (Y_Pos < 10'd195)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd191) && (Y_Pos < 10'd195)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd191) && (Y_Pos < 10'd195)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd191) && (Y_Pos < 10'd195)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd191) && (Y_Pos < 10'd195)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd191) && (Y_Pos < 10'd195)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd191) && (Y_Pos < 10'd195)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd192) && (Y_Pos < 10'd196)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd192) && (Y_Pos < 10'd196)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd192) && (Y_Pos < 10'd196)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd192) && (Y_Pos < 10'd196)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd192) && (Y_Pos < 10'd196)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd192) && (Y_Pos < 10'd196)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd192) && (Y_Pos < 10'd196)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd192) && (Y_Pos < 10'd196)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd193) && (Y_Pos < 10'd197)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd193) && (Y_Pos < 10'd197)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd193) && (Y_Pos < 10'd197)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd193) && (Y_Pos < 10'd197)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd193) && (Y_Pos < 10'd197)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd193) && (Y_Pos < 10'd197)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd193) && (Y_Pos < 10'd197)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd193) && (Y_Pos < 10'd197)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd194) && (Y_Pos < 10'd198)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd194) && (Y_Pos < 10'd198)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd194) && (Y_Pos < 10'd198)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd194) && (Y_Pos < 10'd198)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd194) && (Y_Pos < 10'd198)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd194) && (Y_Pos < 10'd198)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd194) && (Y_Pos < 10'd198)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd194) && (Y_Pos < 10'd198)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd195) && (Y_Pos < 10'd199)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd195) && (Y_Pos < 10'd199)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd195) && (Y_Pos < 10'd199)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd195) && (Y_Pos < 10'd199)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd195) && (Y_Pos < 10'd199)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd195) && (Y_Pos < 10'd199)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd195) && (Y_Pos < 10'd199)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd195) && (Y_Pos < 10'd199)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd196) && (Y_Pos < 10'd200)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd196) && (Y_Pos < 10'd200)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd196) && (Y_Pos < 10'd200)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd196) && (Y_Pos < 10'd200)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd196) && (Y_Pos < 10'd200)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd196) && (Y_Pos < 10'd200)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd196) && (Y_Pos < 10'd200)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd196) && (Y_Pos < 10'd200)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd197) && (Y_Pos < 10'd201)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd197) && (Y_Pos < 10'd201)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd197) && (Y_Pos < 10'd201)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd197) && (Y_Pos < 10'd201)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd197) && (Y_Pos < 10'd201)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd197) && (Y_Pos < 10'd201)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd197) && (Y_Pos < 10'd201)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd197) && (Y_Pos < 10'd201)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd198) && (Y_Pos < 10'd202)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd198) && (Y_Pos < 10'd202)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd198) && (Y_Pos < 10'd202)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd198) && (Y_Pos < 10'd202)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd198) && (Y_Pos < 10'd202)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd198) && (Y_Pos < 10'd202)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd198) && (Y_Pos < 10'd202)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd198) && (Y_Pos < 10'd202)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd199) && (Y_Pos < 10'd203)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd199) && (Y_Pos < 10'd203)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd199) && (Y_Pos < 10'd203)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd199) && (Y_Pos < 10'd203)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd199) && (Y_Pos < 10'd203)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd199) && (Y_Pos < 10'd203)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd199) && (Y_Pos < 10'd203)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd199) && (Y_Pos < 10'd203)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd200) && (Y_Pos < 10'd204)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd200) && (Y_Pos < 10'd204)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd200) && (Y_Pos < 10'd204)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd200) && (Y_Pos < 10'd204)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd200) && (Y_Pos < 10'd204)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd200) && (Y_Pos < 10'd204)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd200) && (Y_Pos < 10'd204)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd200) && (Y_Pos < 10'd204)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd201) && (Y_Pos < 10'd205)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd201) && (Y_Pos < 10'd205)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd201) && (Y_Pos < 10'd205)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd201) && (Y_Pos < 10'd205)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd201) && (Y_Pos < 10'd205)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd201) && (Y_Pos < 10'd205)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd201) && (Y_Pos < 10'd205)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd201) && (Y_Pos < 10'd205)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd202) && (Y_Pos < 10'd206)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd202) && (Y_Pos < 10'd206)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd202) && (Y_Pos < 10'd206)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd202) && (Y_Pos < 10'd206)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd202) && (Y_Pos < 10'd206)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd202) && (Y_Pos < 10'd206)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd202) && (Y_Pos < 10'd206)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd202) && (Y_Pos < 10'd206)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd203) && (Y_Pos < 10'd207)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd203) && (Y_Pos < 10'd207)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd203) && (Y_Pos < 10'd207)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd203) && (Y_Pos < 10'd207)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd203) && (Y_Pos < 10'd207)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd203) && (Y_Pos < 10'd207)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd203) && (Y_Pos < 10'd207)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd203) && (Y_Pos < 10'd207)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd204) && (Y_Pos < 10'd208)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd204) && (Y_Pos < 10'd208)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd204) && (Y_Pos < 10'd208)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd204) && (Y_Pos < 10'd208)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd204) && (Y_Pos < 10'd208)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd204) && (Y_Pos < 10'd208)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd204) && (Y_Pos < 10'd208)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd204) && (Y_Pos < 10'd208)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd205) && (Y_Pos < 10'd209)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd205) && (Y_Pos < 10'd209)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd205) && (Y_Pos < 10'd209)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd205) && (Y_Pos < 10'd209)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd205) && (Y_Pos < 10'd209)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd205) && (Y_Pos < 10'd209)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd205) && (Y_Pos < 10'd209)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd205) && (Y_Pos < 10'd209)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd206) && (Y_Pos < 10'd210)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd206) && (Y_Pos < 10'd210)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd206) && (Y_Pos < 10'd210)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd206) && (Y_Pos < 10'd210)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd206) && (Y_Pos < 10'd210)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd206) && (Y_Pos < 10'd210)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd206) && (Y_Pos < 10'd210)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd206) && (Y_Pos < 10'd210)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd207) && (Y_Pos < 10'd211)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd207) && (Y_Pos < 10'd211)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd207) && (Y_Pos < 10'd211)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd207) && (Y_Pos < 10'd211)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd306) && (Y_Pos > 10'd207) && (Y_Pos < 10'd211)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd333) && (X_Pos < 10'd371) && (Y_Pos > 10'd207) && (Y_Pos < 10'd211)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd207) && (Y_Pos < 10'd211)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd207) && (Y_Pos < 10'd211)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd207) && (Y_Pos < 10'd211)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd207) && (Y_Pos < 10'd211)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd208) && (Y_Pos < 10'd212)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd208) && (Y_Pos < 10'd212)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd208) && (Y_Pos < 10'd212)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd208) && (Y_Pos < 10'd212)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd307) && (Y_Pos > 10'd208) && (Y_Pos < 10'd212)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd332) && (X_Pos < 10'd371) && (Y_Pos > 10'd208) && (Y_Pos < 10'd212)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd208) && (Y_Pos < 10'd212)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd208) && (Y_Pos < 10'd212)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd208) && (Y_Pos < 10'd212)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd208) && (Y_Pos < 10'd212)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd209) && (Y_Pos < 10'd213)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd209) && (Y_Pos < 10'd213)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd209) && (Y_Pos < 10'd213)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd209) && (Y_Pos < 10'd213)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd209) && (Y_Pos < 10'd213)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd302) && (X_Pos < 10'd337) && (Y_Pos > 10'd209) && (Y_Pos < 10'd213)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd209) && (Y_Pos < 10'd213)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd209) && (Y_Pos < 10'd213)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd209) && (Y_Pos < 10'd213)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd209) && (Y_Pos < 10'd213)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd209) && (Y_Pos < 10'd213)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd210) && (Y_Pos < 10'd214)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd210) && (Y_Pos < 10'd214)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd210) && (Y_Pos < 10'd214)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd210) && (Y_Pos < 10'd214)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd210) && (Y_Pos < 10'd214)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd302) && (X_Pos < 10'd337) && (Y_Pos > 10'd210) && (Y_Pos < 10'd214)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd210) && (Y_Pos < 10'd214)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd210) && (Y_Pos < 10'd214)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd210) && (Y_Pos < 10'd214)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd210) && (Y_Pos < 10'd214)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd210) && (Y_Pos < 10'd214)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd211) && (Y_Pos < 10'd215)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd211) && (Y_Pos < 10'd215)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd211) && (Y_Pos < 10'd215)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd211) && (Y_Pos < 10'd215)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd211) && (Y_Pos < 10'd215)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd302) && (X_Pos < 10'd337) && (Y_Pos > 10'd211) && (Y_Pos < 10'd215)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd211) && (Y_Pos < 10'd215)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd211) && (Y_Pos < 10'd215)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd211) && (Y_Pos < 10'd215)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd211) && (Y_Pos < 10'd215)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd211) && (Y_Pos < 10'd215)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd212) && (Y_Pos < 10'd216)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd212) && (Y_Pos < 10'd216)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd212) && (Y_Pos < 10'd216)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd212) && (Y_Pos < 10'd216)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd212) && (Y_Pos < 10'd216)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd274) && (X_Pos < 10'd307) && (Y_Pos > 10'd212) && (Y_Pos < 10'd216)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd332) && (X_Pos < 10'd365) && (Y_Pos > 10'd212) && (Y_Pos < 10'd216)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd212) && (Y_Pos < 10'd216)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd212) && (Y_Pos < 10'd216)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd212) && (Y_Pos < 10'd216)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd212) && (Y_Pos < 10'd216)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd212) && (Y_Pos < 10'd216)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd213) && (Y_Pos < 10'd217)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd213) && (Y_Pos < 10'd217)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd213) && (Y_Pos < 10'd217)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd213) && (Y_Pos < 10'd217)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd213) && (Y_Pos < 10'd217)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd273) && (X_Pos < 10'd306) && (Y_Pos > 10'd213) && (Y_Pos < 10'd217)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd333) && (X_Pos < 10'd366) && (Y_Pos > 10'd213) && (Y_Pos < 10'd217)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd213) && (Y_Pos < 10'd217)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd213) && (Y_Pos < 10'd217)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd213) && (Y_Pos < 10'd217)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd213) && (Y_Pos < 10'd217)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd213) && (Y_Pos < 10'd217)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd192) && (Y_Pos > 10'd214) && (Y_Pos < 10'd218)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd214) && (Y_Pos < 10'd218)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd214) && (Y_Pos < 10'd218)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd214) && (Y_Pos < 10'd218)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd214) && (Y_Pos < 10'd218)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd273) && (X_Pos < 10'd278) && (Y_Pos > 10'd214) && (Y_Pos < 10'd218)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd361) && (X_Pos < 10'd366) && (Y_Pos > 10'd214) && (Y_Pos < 10'd218)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd214) && (Y_Pos < 10'd218)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd214) && (Y_Pos < 10'd218)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd214) && (Y_Pos < 10'd218)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd214) && (Y_Pos < 10'd218)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd447) && (X_Pos < 10'd521) && (Y_Pos > 10'd214) && (Y_Pos < 10'd218)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd188) && (Y_Pos > 10'd215) && (Y_Pos < 10'd219)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd187) && (X_Pos < 10'd192) && (Y_Pos > 10'd215) && (Y_Pos < 10'd219)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd215) && (Y_Pos < 10'd219)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd215) && (Y_Pos < 10'd219)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd215) && (Y_Pos < 10'd219)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd215) && (Y_Pos < 10'd219)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd273) && (X_Pos < 10'd278) && (Y_Pos > 10'd215) && (Y_Pos < 10'd219)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd361) && (X_Pos < 10'd366) && (Y_Pos > 10'd215) && (Y_Pos < 10'd219)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd215) && (Y_Pos < 10'd219)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd215) && (Y_Pos < 10'd219)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd215) && (Y_Pos < 10'd219)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd215) && (Y_Pos < 10'd219)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd447) && (X_Pos < 10'd452) && (Y_Pos > 10'd215) && (Y_Pos < 10'd219)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd451) && (X_Pos < 10'd521) && (Y_Pos > 10'd215) && (Y_Pos < 10'd219)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd216) && (Y_Pos < 10'd220)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd216) && (Y_Pos < 10'd220)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd237) && (X_Pos < 10'd242) && (Y_Pos > 10'd216) && (Y_Pos < 10'd220)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd216) && (Y_Pos < 10'd220)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd273) && (X_Pos < 10'd278) && (Y_Pos > 10'd216) && (Y_Pos < 10'd220)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd361) && (X_Pos < 10'd366) && (Y_Pos > 10'd216) && (Y_Pos < 10'd220)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd216) && (Y_Pos < 10'd220)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd397) && (X_Pos < 10'd402) && (Y_Pos > 10'd216) && (Y_Pos < 10'd220)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd216) && (Y_Pos < 10'd220)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd216) && (Y_Pos < 10'd220)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd193) && (X_Pos < 10'd198) && (Y_Pos > 10'd217) && (Y_Pos < 10'd221)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd227) && (X_Pos < 10'd232) && (Y_Pos > 10'd217) && (Y_Pos < 10'd221)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd236) && (X_Pos < 10'd241) && (Y_Pos > 10'd217) && (Y_Pos < 10'd221)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd217) && (Y_Pos < 10'd221)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd273) && (X_Pos < 10'd278) && (Y_Pos > 10'd217) && (Y_Pos < 10'd221)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd361) && (X_Pos < 10'd366) && (Y_Pos > 10'd217) && (Y_Pos < 10'd221)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd217) && (Y_Pos < 10'd221)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd398) && (X_Pos < 10'd403) && (Y_Pos > 10'd217) && (Y_Pos < 10'd221)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd407) && (X_Pos < 10'd412) && (Y_Pos > 10'd217) && (Y_Pos < 10'd221)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd441) && (X_Pos < 10'd446) && (Y_Pos > 10'd217) && (Y_Pos < 10'd221)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd197) && (Y_Pos > 10'd218) && (Y_Pos < 10'd222)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd227) && (X_Pos < 10'd240) && (Y_Pos > 10'd218) && (Y_Pos < 10'd222)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd218) && (Y_Pos < 10'd222)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd273) && (X_Pos < 10'd278) && (Y_Pos > 10'd218) && (Y_Pos < 10'd222)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd361) && (X_Pos < 10'd366) && (Y_Pos > 10'd218) && (Y_Pos < 10'd222)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd218) && (Y_Pos < 10'd222)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd399) && (X_Pos < 10'd412) && (Y_Pos > 10'd218) && (Y_Pos < 10'd222)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd442) && (X_Pos < 10'd521) && (Y_Pos > 10'd218) && (Y_Pos < 10'd222)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd196) && (Y_Pos > 10'd219) && (Y_Pos < 10'd223)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd229) && (X_Pos < 10'd239) && (Y_Pos > 10'd219) && (Y_Pos < 10'd223)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd219) && (Y_Pos < 10'd223)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd273) && (X_Pos < 10'd278) && (Y_Pos > 10'd219) && (Y_Pos < 10'd223)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd361) && (X_Pos < 10'd366) && (Y_Pos > 10'd219) && (Y_Pos < 10'd223)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd219) && (Y_Pos < 10'd223)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd400) && (X_Pos < 10'd410) && (Y_Pos > 10'd219) && (Y_Pos < 10'd223)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd443) && (X_Pos < 10'd521) && (Y_Pos > 10'd219) && (Y_Pos < 10'd223)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd220) && (Y_Pos < 10'd224)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd273) && (X_Pos < 10'd278) && (Y_Pos > 10'd220) && (Y_Pos < 10'd224)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd361) && (X_Pos < 10'd366) && (Y_Pos > 10'd220) && (Y_Pos < 10'd224)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd220) && (Y_Pos < 10'd224)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd221) && (Y_Pos < 10'd225)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd273) && (X_Pos < 10'd278) && (Y_Pos > 10'd221) && (Y_Pos < 10'd225)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd361) && (X_Pos < 10'd366) && (Y_Pos > 10'd221) && (Y_Pos < 10'd225)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd221) && (Y_Pos < 10'd225)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd222) && (Y_Pos < 10'd226)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd273) && (X_Pos < 10'd278) && (Y_Pos > 10'd222) && (Y_Pos < 10'd226)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd361) && (X_Pos < 10'd366) && (Y_Pos > 10'd222) && (Y_Pos < 10'd226)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd222) && (Y_Pos < 10'd226)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd223) && (Y_Pos < 10'd227)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd273) && (X_Pos < 10'd278) && (Y_Pos > 10'd223) && (Y_Pos < 10'd227)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd361) && (X_Pos < 10'd366) && (Y_Pos > 10'd223) && (Y_Pos < 10'd227)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd223) && (Y_Pos < 10'd227)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd224) && (Y_Pos < 10'd228)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd273) && (X_Pos < 10'd278) && (Y_Pos > 10'd224) && (Y_Pos < 10'd228)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd361) && (X_Pos < 10'd366) && (Y_Pos > 10'd224) && (Y_Pos < 10'd228)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd224) && (Y_Pos < 10'd228)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd225) && (Y_Pos < 10'd229)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd273) && (X_Pos < 10'd278) && (Y_Pos > 10'd225) && (Y_Pos < 10'd229)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd361) && (X_Pos < 10'd366) && (Y_Pos > 10'd225) && (Y_Pos < 10'd229)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd225) && (Y_Pos < 10'd229)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd226) && (Y_Pos < 10'd230)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd273) && (X_Pos < 10'd278) && (Y_Pos > 10'd226) && (Y_Pos < 10'd230)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd361) && (X_Pos < 10'd366) && (Y_Pos > 10'd226) && (Y_Pos < 10'd230)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd226) && (Y_Pos < 10'd230)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd227) && (Y_Pos < 10'd231)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd273) && (X_Pos < 10'd278) && (Y_Pos > 10'd227) && (Y_Pos < 10'd231)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd361) && (X_Pos < 10'd366) && (Y_Pos > 10'd227) && (Y_Pos < 10'd231)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd227) && (Y_Pos < 10'd231)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd228) && (Y_Pos < 10'd232)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd273) && (X_Pos < 10'd278) && (Y_Pos > 10'd228) && (Y_Pos < 10'd232)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd361) && (X_Pos < 10'd366) && (Y_Pos > 10'd228) && (Y_Pos < 10'd232)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd228) && (Y_Pos < 10'd232)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd229) && (Y_Pos < 10'd233)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd273) && (X_Pos < 10'd278) && (Y_Pos > 10'd229) && (Y_Pos < 10'd233)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd361) && (X_Pos < 10'd366) && (Y_Pos > 10'd229) && (Y_Pos < 10'd233)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd229) && (Y_Pos < 10'd233)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd230) && (Y_Pos < 10'd234)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd273) && (X_Pos < 10'd278) && (Y_Pos > 10'd230) && (Y_Pos < 10'd234)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd361) && (X_Pos < 10'd366) && (Y_Pos > 10'd230) && (Y_Pos < 10'd234)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd230) && (Y_Pos < 10'd234)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd231) && (Y_Pos < 10'd235)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd273) && (X_Pos < 10'd278) && (Y_Pos > 10'd231) && (Y_Pos < 10'd235)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd361) && (X_Pos < 10'd366) && (Y_Pos > 10'd231) && (Y_Pos < 10'd235)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd231) && (Y_Pos < 10'd235)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd232) && (Y_Pos < 10'd236)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd273) && (X_Pos < 10'd278) && (Y_Pos > 10'd232) && (Y_Pos < 10'd236)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd361) && (X_Pos < 10'd366) && (Y_Pos > 10'd232) && (Y_Pos < 10'd236)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd232) && (Y_Pos < 10'd236)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd233) && (Y_Pos < 10'd237)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd273) && (X_Pos < 10'd278) && (Y_Pos > 10'd233) && (Y_Pos < 10'd237)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd361) && (X_Pos < 10'd366) && (Y_Pos > 10'd233) && (Y_Pos < 10'd237)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd233) && (Y_Pos < 10'd237)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd234) && (Y_Pos < 10'd238)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd273) && (X_Pos < 10'd278) && (Y_Pos > 10'd234) && (Y_Pos < 10'd238)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd361) && (X_Pos < 10'd366) && (Y_Pos > 10'd234) && (Y_Pos < 10'd238)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd234) && (Y_Pos < 10'd238)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd235) && (Y_Pos < 10'd239)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd273) && (X_Pos < 10'd278) && (Y_Pos > 10'd235) && (Y_Pos < 10'd239)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd361) && (X_Pos < 10'd366) && (Y_Pos > 10'd235) && (Y_Pos < 10'd239)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd235) && (Y_Pos < 10'd239)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd236) && (Y_Pos < 10'd240)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd273) && (X_Pos < 10'd278) && (Y_Pos > 10'd236) && (Y_Pos < 10'd240)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd361) && (X_Pos < 10'd366) && (Y_Pos > 10'd236) && (Y_Pos < 10'd240)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd236) && (Y_Pos < 10'd240)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd237) && (Y_Pos < 10'd241)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd273) && (X_Pos < 10'd278) && (Y_Pos > 10'd237) && (Y_Pos < 10'd241)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd361) && (X_Pos < 10'd366) && (Y_Pos > 10'd237) && (Y_Pos < 10'd241)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd237) && (Y_Pos < 10'd241)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd238) && (Y_Pos < 10'd242)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd273) && (X_Pos < 10'd278) && (Y_Pos > 10'd238) && (Y_Pos < 10'd242)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd361) && (X_Pos < 10'd366) && (Y_Pos > 10'd238) && (Y_Pos < 10'd242)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd238) && (Y_Pos < 10'd242)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd239) && (Y_Pos < 10'd243)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd273) && (X_Pos < 10'd278) && (Y_Pos > 10'd239) && (Y_Pos < 10'd243)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd361) && (X_Pos < 10'd366) && (Y_Pos > 10'd239) && (Y_Pos < 10'd243)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd239) && (Y_Pos < 10'd243)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd240) && (Y_Pos < 10'd244)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd273) && (X_Pos < 10'd278) && (Y_Pos > 10'd240) && (Y_Pos < 10'd244)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd361) && (X_Pos < 10'd366) && (Y_Pos > 10'd240) && (Y_Pos < 10'd244)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd240) && (Y_Pos < 10'd244)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd241) && (Y_Pos < 10'd245)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd273) && (X_Pos < 10'd278) && (Y_Pos > 10'd241) && (Y_Pos < 10'd245)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd361) && (X_Pos < 10'd366) && (Y_Pos > 10'd241) && (Y_Pos < 10'd245)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd241) && (Y_Pos < 10'd245)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd242) && (Y_Pos < 10'd246)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd273) && (X_Pos < 10'd278) && (Y_Pos > 10'd242) && (Y_Pos < 10'd246)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd361) && (X_Pos < 10'd366) && (Y_Pos > 10'd242) && (Y_Pos < 10'd246)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd242) && (Y_Pos < 10'd246)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd243) && (Y_Pos < 10'd247)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd273) && (X_Pos < 10'd278) && (Y_Pos > 10'd243) && (Y_Pos < 10'd247)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd361) && (X_Pos < 10'd366) && (Y_Pos > 10'd243) && (Y_Pos < 10'd247)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd243) && (Y_Pos < 10'd247)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd244) && (Y_Pos < 10'd248)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd273) && (X_Pos < 10'd278) && (Y_Pos > 10'd244) && (Y_Pos < 10'd248)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd361) && (X_Pos < 10'd366) && (Y_Pos > 10'd244) && (Y_Pos < 10'd248)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd244) && (Y_Pos < 10'd248)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd245) && (Y_Pos < 10'd249)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd273) && (X_Pos < 10'd278) && (Y_Pos > 10'd245) && (Y_Pos < 10'd249)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd361) && (X_Pos < 10'd366) && (Y_Pos > 10'd245) && (Y_Pos < 10'd249)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd245) && (Y_Pos < 10'd249)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd196) && (Y_Pos > 10'd246) && (Y_Pos < 10'd250)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd229) && (X_Pos < 10'd239) && (Y_Pos > 10'd246) && (Y_Pos < 10'd250)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd246) && (Y_Pos < 10'd250)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd273) && (X_Pos < 10'd278) && (Y_Pos > 10'd246) && (Y_Pos < 10'd250)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd361) && (X_Pos < 10'd366) && (Y_Pos > 10'd246) && (Y_Pos < 10'd250)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd246) && (Y_Pos < 10'd250)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd400) && (X_Pos < 10'd410) && (Y_Pos > 10'd246) && (Y_Pos < 10'd250)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd443) && (X_Pos < 10'd521) && (Y_Pos > 10'd246) && (Y_Pos < 10'd250)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd197) && (Y_Pos > 10'd247) && (Y_Pos < 10'd251)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd228) && (X_Pos < 10'd240) && (Y_Pos > 10'd247) && (Y_Pos < 10'd251)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd247) && (Y_Pos < 10'd251)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd273) && (X_Pos < 10'd278) && (Y_Pos > 10'd247) && (Y_Pos < 10'd251)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd361) && (X_Pos < 10'd366) && (Y_Pos > 10'd247) && (Y_Pos < 10'd251)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd247) && (Y_Pos < 10'd251)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd399) && (X_Pos < 10'd411) && (Y_Pos > 10'd247) && (Y_Pos < 10'd251)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd442) && (X_Pos < 10'd521) && (Y_Pos > 10'd247) && (Y_Pos < 10'd251)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd193) && (X_Pos < 10'd198) && (Y_Pos > 10'd248) && (Y_Pos < 10'd252)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd227) && (X_Pos < 10'd232) && (Y_Pos > 10'd248) && (Y_Pos < 10'd252)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd236) && (X_Pos < 10'd241) && (Y_Pos > 10'd248) && (Y_Pos < 10'd252)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd248) && (Y_Pos < 10'd252)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd273) && (X_Pos < 10'd278) && (Y_Pos > 10'd248) && (Y_Pos < 10'd252)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd361) && (X_Pos < 10'd366) && (Y_Pos > 10'd248) && (Y_Pos < 10'd252)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd248) && (Y_Pos < 10'd252)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd398) && (X_Pos < 10'd403) && (Y_Pos > 10'd248) && (Y_Pos < 10'd252)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd407) && (X_Pos < 10'd412) && (Y_Pos > 10'd248) && (Y_Pos < 10'd252)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd441) && (X_Pos < 10'd446) && (Y_Pos > 10'd248) && (Y_Pos < 10'd252)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd194) && (X_Pos < 10'd199) && (Y_Pos > 10'd249) && (Y_Pos < 10'd253)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd249) && (Y_Pos < 10'd253)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd237) && (X_Pos < 10'd242) && (Y_Pos > 10'd249) && (Y_Pos < 10'd253)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd249) && (Y_Pos < 10'd253)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd273) && (X_Pos < 10'd278) && (Y_Pos > 10'd249) && (Y_Pos < 10'd253)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd361) && (X_Pos < 10'd366) && (Y_Pos > 10'd249) && (Y_Pos < 10'd253)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd249) && (Y_Pos < 10'd253)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd397) && (X_Pos < 10'd402) && (Y_Pos > 10'd249) && (Y_Pos < 10'd253)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd249) && (Y_Pos < 10'd253)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd440) && (X_Pos < 10'd445) && (Y_Pos > 10'd249) && (Y_Pos < 10'd253)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd250) && (Y_Pos < 10'd254)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd250) && (Y_Pos < 10'd254)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd250) && (Y_Pos < 10'd254)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd250) && (Y_Pos < 10'd254)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd273) && (X_Pos < 10'd278) && (Y_Pos > 10'd250) && (Y_Pos < 10'd254)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd361) && (X_Pos < 10'd366) && (Y_Pos > 10'd250) && (Y_Pos < 10'd254)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd250) && (Y_Pos < 10'd254)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd250) && (Y_Pos < 10'd254)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd250) && (Y_Pos < 10'd254)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd250) && (Y_Pos < 10'd254)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd192) && (Y_Pos > 10'd251) && (Y_Pos < 10'd255)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd251) && (Y_Pos < 10'd255)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd251) && (Y_Pos < 10'd255)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd251) && (Y_Pos < 10'd255)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd251) && (Y_Pos < 10'd255)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd273) && (X_Pos < 10'd278) && (Y_Pos > 10'd251) && (Y_Pos < 10'd255)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd361) && (X_Pos < 10'd366) && (Y_Pos > 10'd251) && (Y_Pos < 10'd255)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd251) && (Y_Pos < 10'd255)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd251) && (Y_Pos < 10'd255)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd251) && (Y_Pos < 10'd255)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd251) && (Y_Pos < 10'd255)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd447) && (X_Pos < 10'd521) && (Y_Pos > 10'd251) && (Y_Pos < 10'd255)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd194) && (Y_Pos > 10'd252) && (Y_Pos < 10'd256)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd252) && (Y_Pos < 10'd256)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd252) && (Y_Pos < 10'd256)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd252) && (Y_Pos < 10'd256)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd252) && (Y_Pos < 10'd256)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd273) && (X_Pos < 10'd366) && (Y_Pos > 10'd252) && (Y_Pos < 10'd256)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd252) && (Y_Pos < 10'd256)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd252) && (Y_Pos < 10'd256)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd252) && (Y_Pos < 10'd256)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd252) && (Y_Pos < 10'd256)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd521) && (Y_Pos > 10'd252) && (Y_Pos < 10'd256)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd253) && (Y_Pos < 10'd257)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd253) && (Y_Pos < 10'd257)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd253) && (Y_Pos < 10'd257)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd253) && (Y_Pos < 10'd257)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd253) && (Y_Pos < 10'd257)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd273) && (X_Pos < 10'd366) && (Y_Pos > 10'd253) && (Y_Pos < 10'd257)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd253) && (Y_Pos < 10'd257)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd253) && (Y_Pos < 10'd257)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd253) && (Y_Pos < 10'd257)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd253) && (Y_Pos < 10'd257)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd253) && (Y_Pos < 10'd257)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd254) && (Y_Pos < 10'd258)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd254) && (Y_Pos < 10'd258)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd254) && (Y_Pos < 10'd258)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd254) && (Y_Pos < 10'd258)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd254) && (Y_Pos < 10'd258)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd254) && (Y_Pos < 10'd258)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd254) && (Y_Pos < 10'd258)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd254) && (Y_Pos < 10'd258)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd254) && (Y_Pos < 10'd258)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd254) && (Y_Pos < 10'd258)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd255) && (Y_Pos < 10'd259)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd255) && (Y_Pos < 10'd259)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd255) && (Y_Pos < 10'd259)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd255) && (Y_Pos < 10'd259)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd255) && (Y_Pos < 10'd259)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd255) && (Y_Pos < 10'd259)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd255) && (Y_Pos < 10'd259)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd255) && (Y_Pos < 10'd259)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd255) && (Y_Pos < 10'd259)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd255) && (Y_Pos < 10'd259)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd256) && (Y_Pos < 10'd260)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd256) && (Y_Pos < 10'd260)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd256) && (Y_Pos < 10'd260)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd256) && (Y_Pos < 10'd260)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd256) && (Y_Pos < 10'd260)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd256) && (Y_Pos < 10'd260)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd256) && (Y_Pos < 10'd260)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd256) && (Y_Pos < 10'd260)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd256) && (Y_Pos < 10'd260)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd256) && (Y_Pos < 10'd260)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd257) && (Y_Pos < 10'd261)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd257) && (Y_Pos < 10'd261)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd257) && (Y_Pos < 10'd261)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd257) && (Y_Pos < 10'd261)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd371) && (Y_Pos > 10'd257) && (Y_Pos < 10'd261)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd257) && (Y_Pos < 10'd261)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd257) && (Y_Pos < 10'd261)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd257) && (Y_Pos < 10'd261)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd257) && (Y_Pos < 10'd261)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd258) && (Y_Pos < 10'd262)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd258) && (Y_Pos < 10'd262)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd258) && (Y_Pos < 10'd262)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd258) && (Y_Pos < 10'd262)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd371) && (Y_Pos > 10'd258) && (Y_Pos < 10'd262)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd258) && (Y_Pos < 10'd262)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd258) && (Y_Pos < 10'd262)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd258) && (Y_Pos < 10'd262)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd258) && (Y_Pos < 10'd262)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd259) && (Y_Pos < 10'd263)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd259) && (Y_Pos < 10'd263)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd259) && (Y_Pos < 10'd263)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd259) && (Y_Pos < 10'd263)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd259) && (Y_Pos < 10'd263)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd259) && (Y_Pos < 10'd263)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd259) && (Y_Pos < 10'd263)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd259) && (Y_Pos < 10'd263)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd260) && (Y_Pos < 10'd264)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd260) && (Y_Pos < 10'd264)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd260) && (Y_Pos < 10'd264)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd260) && (Y_Pos < 10'd264)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd260) && (Y_Pos < 10'd264)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd260) && (Y_Pos < 10'd264)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd260) && (Y_Pos < 10'd264)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd260) && (Y_Pos < 10'd264)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd261) && (Y_Pos < 10'd265)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd261) && (Y_Pos < 10'd265)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd261) && (Y_Pos < 10'd265)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd261) && (Y_Pos < 10'd265)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd261) && (Y_Pos < 10'd265)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd261) && (Y_Pos < 10'd265)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd261) && (Y_Pos < 10'd265)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd261) && (Y_Pos < 10'd265)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd262) && (Y_Pos < 10'd266)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd262) && (Y_Pos < 10'd266)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd262) && (Y_Pos < 10'd266)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd262) && (Y_Pos < 10'd266)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd262) && (Y_Pos < 10'd266)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd262) && (Y_Pos < 10'd266)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd262) && (Y_Pos < 10'd266)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd262) && (Y_Pos < 10'd266)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd263) && (Y_Pos < 10'd267)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd263) && (Y_Pos < 10'd267)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd263) && (Y_Pos < 10'd267)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd263) && (Y_Pos < 10'd267)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd263) && (Y_Pos < 10'd267)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd263) && (Y_Pos < 10'd267)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd263) && (Y_Pos < 10'd267)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd263) && (Y_Pos < 10'd267)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd264) && (Y_Pos < 10'd268)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd264) && (Y_Pos < 10'd268)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd264) && (Y_Pos < 10'd268)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd264) && (Y_Pos < 10'd268)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd264) && (Y_Pos < 10'd268)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd264) && (Y_Pos < 10'd268)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd264) && (Y_Pos < 10'd268)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd264) && (Y_Pos < 10'd268)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd265) && (Y_Pos < 10'd269)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd265) && (Y_Pos < 10'd269)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd265) && (Y_Pos < 10'd269)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd265) && (Y_Pos < 10'd269)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd265) && (Y_Pos < 10'd269)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd265) && (Y_Pos < 10'd269)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd265) && (Y_Pos < 10'd269)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd265) && (Y_Pos < 10'd269)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd266) && (Y_Pos < 10'd270)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd266) && (Y_Pos < 10'd270)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd266) && (Y_Pos < 10'd270)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd266) && (Y_Pos < 10'd270)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd266) && (Y_Pos < 10'd270)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd266) && (Y_Pos < 10'd270)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd266) && (Y_Pos < 10'd270)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd266) && (Y_Pos < 10'd270)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd267) && (Y_Pos < 10'd271)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd267) && (Y_Pos < 10'd271)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd267) && (Y_Pos < 10'd271)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd267) && (Y_Pos < 10'd271)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd267) && (Y_Pos < 10'd271)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd267) && (Y_Pos < 10'd271)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd267) && (Y_Pos < 10'd271)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd267) && (Y_Pos < 10'd271)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd268) && (Y_Pos < 10'd272)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd268) && (Y_Pos < 10'd272)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd268) && (Y_Pos < 10'd272)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd268) && (Y_Pos < 10'd272)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd268) && (Y_Pos < 10'd272)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd268) && (Y_Pos < 10'd272)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd268) && (Y_Pos < 10'd272)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd268) && (Y_Pos < 10'd272)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd269) && (Y_Pos < 10'd273)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd269) && (Y_Pos < 10'd273)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd269) && (Y_Pos < 10'd273)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd269) && (Y_Pos < 10'd273)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd269) && (Y_Pos < 10'd273)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd269) && (Y_Pos < 10'd273)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd269) && (Y_Pos < 10'd273)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd269) && (Y_Pos < 10'd273)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd270) && (Y_Pos < 10'd274)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd270) && (Y_Pos < 10'd274)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd270) && (Y_Pos < 10'd274)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd270) && (Y_Pos < 10'd274)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd270) && (Y_Pos < 10'd274)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd270) && (Y_Pos < 10'd274)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd270) && (Y_Pos < 10'd274)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd270) && (Y_Pos < 10'd274)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd271) && (Y_Pos < 10'd275)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd271) && (Y_Pos < 10'd275)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd271) && (Y_Pos < 10'd275)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd271) && (Y_Pos < 10'd275)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd271) && (Y_Pos < 10'd275)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd271) && (Y_Pos < 10'd275)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd271) && (Y_Pos < 10'd275)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd271) && (Y_Pos < 10'd275)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd272) && (Y_Pos < 10'd276)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd272) && (Y_Pos < 10'd276)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd272) && (Y_Pos < 10'd276)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd272) && (Y_Pos < 10'd276)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd272) && (Y_Pos < 10'd276)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd272) && (Y_Pos < 10'd276)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd272) && (Y_Pos < 10'd276)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd272) && (Y_Pos < 10'd276)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd273) && (Y_Pos < 10'd277)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd273) && (Y_Pos < 10'd277)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd273) && (Y_Pos < 10'd277)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd273) && (Y_Pos < 10'd277)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd273) && (Y_Pos < 10'd277)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd273) && (Y_Pos < 10'd277)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd273) && (Y_Pos < 10'd277)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd273) && (Y_Pos < 10'd277)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd274) && (Y_Pos < 10'd278)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd274) && (Y_Pos < 10'd278)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd274) && (Y_Pos < 10'd278)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd274) && (Y_Pos < 10'd278)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd274) && (Y_Pos < 10'd278)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd274) && (Y_Pos < 10'd278)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd274) && (Y_Pos < 10'd278)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd274) && (Y_Pos < 10'd278)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd275) && (Y_Pos < 10'd279)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd275) && (Y_Pos < 10'd279)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd275) && (Y_Pos < 10'd279)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd275) && (Y_Pos < 10'd279)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd275) && (Y_Pos < 10'd279)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd275) && (Y_Pos < 10'd279)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd275) && (Y_Pos < 10'd279)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd275) && (Y_Pos < 10'd279)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd276) && (Y_Pos < 10'd280)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd276) && (Y_Pos < 10'd280)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd276) && (Y_Pos < 10'd280)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd276) && (Y_Pos < 10'd280)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd276) && (Y_Pos < 10'd280)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd276) && (Y_Pos < 10'd280)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd276) && (Y_Pos < 10'd280)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd276) && (Y_Pos < 10'd280)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd277) && (Y_Pos < 10'd281)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd277) && (Y_Pos < 10'd281)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd277) && (Y_Pos < 10'd281)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd277) && (Y_Pos < 10'd281)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd277) && (Y_Pos < 10'd281)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd277) && (Y_Pos < 10'd281)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd277) && (Y_Pos < 10'd281)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd277) && (Y_Pos < 10'd281)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd278) && (Y_Pos < 10'd282)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd278) && (Y_Pos < 10'd282)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd278) && (Y_Pos < 10'd282)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd278) && (Y_Pos < 10'd282)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd278) && (Y_Pos < 10'd282)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd278) && (Y_Pos < 10'd282)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd278) && (Y_Pos < 10'd282)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd278) && (Y_Pos < 10'd282)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd279) && (Y_Pos < 10'd283)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd279) && (Y_Pos < 10'd283)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd279) && (Y_Pos < 10'd283)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd279) && (Y_Pos < 10'd283)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd279) && (Y_Pos < 10'd283)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd279) && (Y_Pos < 10'd283)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd279) && (Y_Pos < 10'd283)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd279) && (Y_Pos < 10'd283)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd280) && (Y_Pos < 10'd284)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd280) && (Y_Pos < 10'd284)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd280) && (Y_Pos < 10'd284)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd280) && (Y_Pos < 10'd284)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd280) && (Y_Pos < 10'd284)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd280) && (Y_Pos < 10'd284)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd280) && (Y_Pos < 10'd284)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd280) && (Y_Pos < 10'd284)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd281) && (Y_Pos < 10'd285)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd281) && (Y_Pos < 10'd285)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd281) && (Y_Pos < 10'd285)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd281) && (Y_Pos < 10'd285)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd281) && (Y_Pos < 10'd285)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd281) && (Y_Pos < 10'd285)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd281) && (Y_Pos < 10'd285)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd281) && (Y_Pos < 10'd285)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd282) && (Y_Pos < 10'd286)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd282) && (Y_Pos < 10'd286)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd282) && (Y_Pos < 10'd286)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd282) && (Y_Pos < 10'd286)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd282) && (Y_Pos < 10'd286)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd282) && (Y_Pos < 10'd286)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd282) && (Y_Pos < 10'd286)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd282) && (Y_Pos < 10'd286)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd283) && (Y_Pos < 10'd287)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd283) && (Y_Pos < 10'd287)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd283) && (Y_Pos < 10'd287)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd283) && (Y_Pos < 10'd287)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd283) && (Y_Pos < 10'd287)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd283) && (Y_Pos < 10'd287)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd283) && (Y_Pos < 10'd287)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd283) && (Y_Pos < 10'd287)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd284) && (Y_Pos < 10'd288)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd284) && (Y_Pos < 10'd288)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd284) && (Y_Pos < 10'd288)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd284) && (Y_Pos < 10'd288)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd284) && (Y_Pos < 10'd288)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd284) && (Y_Pos < 10'd288)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd284) && (Y_Pos < 10'd288)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd284) && (Y_Pos < 10'd288)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd285) && (Y_Pos < 10'd289)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd285) && (Y_Pos < 10'd289)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd285) && (Y_Pos < 10'd289)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd285) && (Y_Pos < 10'd289)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd272) && (X_Pos < 10'd367) && (Y_Pos > 10'd285) && (Y_Pos < 10'd289)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd285) && (Y_Pos < 10'd289)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd285) && (Y_Pos < 10'd289)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd285) && (Y_Pos < 10'd289)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd285) && (Y_Pos < 10'd289)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd286) && (Y_Pos < 10'd290)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd286) && (Y_Pos < 10'd290)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd286) && (Y_Pos < 10'd290)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd286) && (Y_Pos < 10'd290)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd270) && (X_Pos < 10'd275) && (Y_Pos > 10'd286) && (Y_Pos < 10'd290)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd364) && (X_Pos < 10'd369) && (Y_Pos > 10'd286) && (Y_Pos < 10'd290)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd286) && (Y_Pos < 10'd290)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd286) && (Y_Pos < 10'd290)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd286) && (Y_Pos < 10'd290)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd286) && (Y_Pos < 10'd290)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd287) && (Y_Pos < 10'd291)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd287) && (Y_Pos < 10'd291)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd287) && (Y_Pos < 10'd291)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd287) && (Y_Pos < 10'd291)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd270) && (X_Pos < 10'd275) && (Y_Pos > 10'd287) && (Y_Pos < 10'd291)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd364) && (X_Pos < 10'd369) && (Y_Pos > 10'd287) && (Y_Pos < 10'd291)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd287) && (Y_Pos < 10'd291)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd287) && (Y_Pos < 10'd291)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd287) && (Y_Pos < 10'd291)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd287) && (Y_Pos < 10'd291)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd288) && (Y_Pos < 10'd292)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd288) && (Y_Pos < 10'd292)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd288) && (Y_Pos < 10'd292)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd288) && (Y_Pos < 10'd292)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd288) && (Y_Pos < 10'd292)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd288) && (Y_Pos < 10'd292)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd288) && (Y_Pos < 10'd292)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd288) && (Y_Pos < 10'd292)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd288) && (Y_Pos < 10'd292)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd288) && (Y_Pos < 10'd292)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd289) && (Y_Pos < 10'd293)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd289) && (Y_Pos < 10'd293)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd289) && (Y_Pos < 10'd293)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd289) && (Y_Pos < 10'd293)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd289) && (Y_Pos < 10'd293)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd289) && (Y_Pos < 10'd293)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd289) && (Y_Pos < 10'd293)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd289) && (Y_Pos < 10'd293)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd289) && (Y_Pos < 10'd293)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd289) && (Y_Pos < 10'd293)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd194) && (Y_Pos > 10'd290) && (Y_Pos < 10'd294)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd290) && (Y_Pos < 10'd294)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd290) && (Y_Pos < 10'd294)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd290) && (Y_Pos < 10'd294)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd290) && (Y_Pos < 10'd294)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd290) && (Y_Pos < 10'd294)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd290) && (Y_Pos < 10'd294)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd290) && (Y_Pos < 10'd294)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd290) && (Y_Pos < 10'd294)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd450) && (Y_Pos > 10'd290) && (Y_Pos < 10'd294)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd125) && (X_Pos < 10'd193) && (Y_Pos > 10'd291) && (Y_Pos < 10'd295)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd291) && (Y_Pos < 10'd295)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd291) && (Y_Pos < 10'd295)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd291) && (Y_Pos < 10'd295)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd291) && (Y_Pos < 10'd295)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd291) && (Y_Pos < 10'd295)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd291) && (Y_Pos < 10'd295)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd291) && (Y_Pos < 10'd295)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd291) && (Y_Pos < 10'd295)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd446) && (X_Pos < 10'd514) && (Y_Pos > 10'd291) && (Y_Pos < 10'd295)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd125) && (X_Pos < 10'd192) && (Y_Pos > 10'd292) && (Y_Pos < 10'd296)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd292) && (Y_Pos < 10'd296)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd292) && (Y_Pos < 10'd296)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd292) && (Y_Pos < 10'd296)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd292) && (Y_Pos < 10'd296)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd292) && (Y_Pos < 10'd296)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd292) && (Y_Pos < 10'd296)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd292) && (Y_Pos < 10'd296)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd292) && (Y_Pos < 10'd296)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd447) && (X_Pos < 10'd514) && (Y_Pos > 10'd292) && (Y_Pos < 10'd296)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd122) && (X_Pos < 10'd128) && (Y_Pos > 10'd293) && (Y_Pos < 10'd297)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd293) && (Y_Pos < 10'd297)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd293) && (Y_Pos < 10'd297)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd293) && (Y_Pos < 10'd297)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd293) && (Y_Pos < 10'd297)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd293) && (Y_Pos < 10'd297)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd293) && (Y_Pos < 10'd297)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd293) && (Y_Pos < 10'd297)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd293) && (Y_Pos < 10'd297)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd517) && (Y_Pos > 10'd293) && (Y_Pos < 10'd297)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd120) && (X_Pos < 10'd127) && (Y_Pos > 10'd294) && (Y_Pos < 10'd298)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd193) && (X_Pos < 10'd198) && (Y_Pos > 10'd294) && (Y_Pos < 10'd298)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd226) && (X_Pos < 10'd231) && (Y_Pos > 10'd294) && (Y_Pos < 10'd298)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd236) && (X_Pos < 10'd241) && (Y_Pos > 10'd294) && (Y_Pos < 10'd298)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd269) && (X_Pos < 10'd274) && (Y_Pos > 10'd294) && (Y_Pos < 10'd298)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd365) && (X_Pos < 10'd370) && (Y_Pos > 10'd294) && (Y_Pos < 10'd298)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd398) && (X_Pos < 10'd403) && (Y_Pos > 10'd294) && (Y_Pos < 10'd298)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd408) && (X_Pos < 10'd413) && (Y_Pos > 10'd294) && (Y_Pos < 10'd298)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd441) && (X_Pos < 10'd446) && (Y_Pos > 10'd294) && (Y_Pos < 10'd298)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd512) && (X_Pos < 10'd519) && (Y_Pos > 10'd294) && (Y_Pos < 10'd298)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd120) && (X_Pos < 10'd125) && (Y_Pos > 10'd295) && (Y_Pos < 10'd299)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd193) && (X_Pos < 10'd198) && (Y_Pos > 10'd295) && (Y_Pos < 10'd299)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd227) && (X_Pos < 10'd232) && (Y_Pos > 10'd295) && (Y_Pos < 10'd299)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd236) && (X_Pos < 10'd241) && (Y_Pos > 10'd295) && (Y_Pos < 10'd299)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd270) && (X_Pos < 10'd275) && (Y_Pos > 10'd295) && (Y_Pos < 10'd299)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd364) && (X_Pos < 10'd369) && (Y_Pos > 10'd295) && (Y_Pos < 10'd299)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd398) && (X_Pos < 10'd403) && (Y_Pos > 10'd295) && (Y_Pos < 10'd299)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd407) && (X_Pos < 10'd412) && (Y_Pos > 10'd295) && (Y_Pos < 10'd299)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd441) && (X_Pos < 10'd446) && (Y_Pos > 10'd295) && (Y_Pos < 10'd299)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd514) && (X_Pos < 10'd519) && (Y_Pos > 10'd295) && (Y_Pos < 10'd299)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd120) && (X_Pos < 10'd125) && (Y_Pos > 10'd296) && (Y_Pos < 10'd300)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd127) && (X_Pos < 10'd196) && (Y_Pos > 10'd296) && (Y_Pos < 10'd300)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd229) && (X_Pos < 10'd239) && (Y_Pos > 10'd296) && (Y_Pos < 10'd300)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd271) && (X_Pos < 10'd312) && (Y_Pos > 10'd296) && (Y_Pos < 10'd300)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd327) && (X_Pos < 10'd368) && (Y_Pos > 10'd296) && (Y_Pos < 10'd300)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd400) && (X_Pos < 10'd410) && (Y_Pos > 10'd296) && (Y_Pos < 10'd300)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd443) && (X_Pos < 10'd512) && (Y_Pos > 10'd296) && (Y_Pos < 10'd300)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd514) && (X_Pos < 10'd519) && (Y_Pos > 10'd296) && (Y_Pos < 10'd300)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd120) && (X_Pos < 10'd124) && (Y_Pos > 10'd297) && (Y_Pos < 10'd301)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd126) && (X_Pos < 10'd196) && (Y_Pos > 10'd297) && (Y_Pos < 10'd301)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd229) && (X_Pos < 10'd238) && (Y_Pos > 10'd297) && (Y_Pos < 10'd301)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd272) && (X_Pos < 10'd313) && (Y_Pos > 10'd297) && (Y_Pos < 10'd301)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd326) && (X_Pos < 10'd367) && (Y_Pos > 10'd297) && (Y_Pos < 10'd301)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd401) && (X_Pos < 10'd410) && (Y_Pos > 10'd297) && (Y_Pos < 10'd301)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd443) && (X_Pos < 10'd513) && (Y_Pos > 10'd297) && (Y_Pos < 10'd301)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd515) && (X_Pos < 10'd519) && (Y_Pos > 10'd297) && (Y_Pos < 10'd301)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd298) && (Y_Pos < 10'd302)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd125) && (X_Pos < 10'd130) && (Y_Pos > 10'd298) && (Y_Pos < 10'd302)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd309) && (X_Pos < 10'd314) && (Y_Pos > 10'd298) && (Y_Pos < 10'd302)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd325) && (X_Pos < 10'd330) && (Y_Pos > 10'd298) && (Y_Pos < 10'd302)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd509) && (X_Pos < 10'd514) && (Y_Pos > 10'd298) && (Y_Pos < 10'd302)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd298) && (Y_Pos < 10'd302)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd299) && (Y_Pos < 10'd303)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd129) && (Y_Pos > 10'd299) && (Y_Pos < 10'd303)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd310) && (X_Pos < 10'd315) && (Y_Pos > 10'd299) && (Y_Pos < 10'd303)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd324) && (X_Pos < 10'd329) && (Y_Pos > 10'd299) && (Y_Pos < 10'd303)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd510) && (X_Pos < 10'd516) && (Y_Pos > 10'd299) && (Y_Pos < 10'd303)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd299) && (Y_Pos < 10'd303)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd300) && (Y_Pos < 10'd304)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd300) && (Y_Pos < 10'd304)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd300) && (Y_Pos < 10'd304)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd300) && (Y_Pos < 10'd304)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd300) && (Y_Pos < 10'd304)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd300) && (Y_Pos < 10'd304)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd301) && (Y_Pos < 10'd305)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd301) && (Y_Pos < 10'd305)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd301) && (Y_Pos < 10'd305)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd301) && (Y_Pos < 10'd305)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd301) && (Y_Pos < 10'd305)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd301) && (Y_Pos < 10'd305)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd302) && (Y_Pos < 10'd306)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd302) && (Y_Pos < 10'd306)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd302) && (Y_Pos < 10'd306)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd302) && (Y_Pos < 10'd306)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd302) && (Y_Pos < 10'd306)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd302) && (Y_Pos < 10'd306)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd303) && (Y_Pos < 10'd307)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd303) && (Y_Pos < 10'd307)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd303) && (Y_Pos < 10'd307)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd303) && (Y_Pos < 10'd307)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd303) && (Y_Pos < 10'd307)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd303) && (Y_Pos < 10'd307)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd304) && (Y_Pos < 10'd308)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd304) && (Y_Pos < 10'd308)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd304) && (Y_Pos < 10'd308)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd304) && (Y_Pos < 10'd308)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd304) && (Y_Pos < 10'd308)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd304) && (Y_Pos < 10'd308)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd305) && (Y_Pos < 10'd309)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd305) && (Y_Pos < 10'd309)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd305) && (Y_Pos < 10'd309)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd305) && (Y_Pos < 10'd309)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd305) && (Y_Pos < 10'd309)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd305) && (Y_Pos < 10'd309)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd306) && (Y_Pos < 10'd310)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd306) && (Y_Pos < 10'd310)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd306) && (Y_Pos < 10'd310)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd306) && (Y_Pos < 10'd310)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd306) && (Y_Pos < 10'd310)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd306) && (Y_Pos < 10'd310)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd307) && (Y_Pos < 10'd311)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd307) && (Y_Pos < 10'd311)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd307) && (Y_Pos < 10'd311)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd307) && (Y_Pos < 10'd311)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd307) && (Y_Pos < 10'd311)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd307) && (Y_Pos < 10'd311)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd308) && (Y_Pos < 10'd312)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd308) && (Y_Pos < 10'd312)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd308) && (Y_Pos < 10'd312)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd308) && (Y_Pos < 10'd312)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd308) && (Y_Pos < 10'd312)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd308) && (Y_Pos < 10'd312)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd309) && (Y_Pos < 10'd313)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd309) && (Y_Pos < 10'd313)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd309) && (Y_Pos < 10'd313)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd309) && (Y_Pos < 10'd313)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd309) && (Y_Pos < 10'd313)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd309) && (Y_Pos < 10'd313)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd310) && (Y_Pos < 10'd314)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd310) && (Y_Pos < 10'd314)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd310) && (Y_Pos < 10'd314)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd310) && (Y_Pos < 10'd314)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd310) && (Y_Pos < 10'd314)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd310) && (Y_Pos < 10'd314)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd311) && (Y_Pos < 10'd315)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd311) && (Y_Pos < 10'd315)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd311) && (Y_Pos < 10'd315)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd311) && (Y_Pos < 10'd315)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd311) && (Y_Pos < 10'd315)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd311) && (Y_Pos < 10'd315)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd312) && (Y_Pos < 10'd316)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd312) && (Y_Pos < 10'd316)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd312) && (Y_Pos < 10'd316)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd312) && (Y_Pos < 10'd316)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd312) && (Y_Pos < 10'd316)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd312) && (Y_Pos < 10'd316)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd313) && (Y_Pos < 10'd317)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd313) && (Y_Pos < 10'd317)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd313) && (Y_Pos < 10'd317)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd313) && (Y_Pos < 10'd317)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd313) && (Y_Pos < 10'd317)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd313) && (Y_Pos < 10'd317)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd314) && (Y_Pos < 10'd318)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd314) && (Y_Pos < 10'd318)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd314) && (Y_Pos < 10'd318)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd314) && (Y_Pos < 10'd318)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd314) && (Y_Pos < 10'd318)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd314) && (Y_Pos < 10'd318)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd315) && (Y_Pos < 10'd319)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd315) && (Y_Pos < 10'd319)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd315) && (Y_Pos < 10'd319)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd315) && (Y_Pos < 10'd319)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd315) && (Y_Pos < 10'd319)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd315) && (Y_Pos < 10'd319)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd316) && (Y_Pos < 10'd320)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd316) && (Y_Pos < 10'd320)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd316) && (Y_Pos < 10'd320)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd316) && (Y_Pos < 10'd320)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd316) && (Y_Pos < 10'd320)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd316) && (Y_Pos < 10'd320)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd317) && (Y_Pos < 10'd321)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd317) && (Y_Pos < 10'd321)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd317) && (Y_Pos < 10'd321)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd317) && (Y_Pos < 10'd321)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd317) && (Y_Pos < 10'd321)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd317) && (Y_Pos < 10'd321)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd318) && (Y_Pos < 10'd322)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd318) && (Y_Pos < 10'd322)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd318) && (Y_Pos < 10'd322)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd318) && (Y_Pos < 10'd322)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd318) && (Y_Pos < 10'd322)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd318) && (Y_Pos < 10'd322)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd319) && (Y_Pos < 10'd323)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd319) && (Y_Pos < 10'd323)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd319) && (Y_Pos < 10'd323)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd319) && (Y_Pos < 10'd323)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd319) && (Y_Pos < 10'd323)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd319) && (Y_Pos < 10'd323)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd320) && (Y_Pos < 10'd324)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd320) && (Y_Pos < 10'd324)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd320) && (Y_Pos < 10'd324)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd320) && (Y_Pos < 10'd324)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd320) && (Y_Pos < 10'd324)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd320) && (Y_Pos < 10'd324)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd321) && (Y_Pos < 10'd325)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd321) && (Y_Pos < 10'd325)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd321) && (Y_Pos < 10'd325)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd321) && (Y_Pos < 10'd325)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd321) && (Y_Pos < 10'd325)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd321) && (Y_Pos < 10'd325)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd322) && (Y_Pos < 10'd326)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd322) && (Y_Pos < 10'd326)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd322) && (Y_Pos < 10'd326)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd322) && (Y_Pos < 10'd326)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd322) && (Y_Pos < 10'd326)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd322) && (Y_Pos < 10'd326)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd323) && (Y_Pos < 10'd327)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd323) && (Y_Pos < 10'd327)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd158) && (X_Pos < 10'd196) && (Y_Pos > 10'd323) && (Y_Pos < 10'd327)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd229) && (X_Pos < 10'd281) && (Y_Pos > 10'd323) && (Y_Pos < 10'd327)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd323) && (Y_Pos < 10'd327)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd323) && (Y_Pos < 10'd327)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd358) && (X_Pos < 10'd410) && (Y_Pos > 10'd323) && (Y_Pos < 10'd327)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd443) && (X_Pos < 10'd481) && (Y_Pos > 10'd323) && (Y_Pos < 10'd327)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd323) && (Y_Pos < 10'd327)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd323) && (Y_Pos < 10'd327)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd324) && (Y_Pos < 10'd328)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd324) && (Y_Pos < 10'd328)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd157) && (X_Pos < 10'd196) && (Y_Pos > 10'd324) && (Y_Pos < 10'd328)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd229) && (X_Pos < 10'd282) && (Y_Pos > 10'd324) && (Y_Pos < 10'd328)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd324) && (Y_Pos < 10'd328)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd324) && (Y_Pos < 10'd328)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd357) && (X_Pos < 10'd410) && (Y_Pos > 10'd324) && (Y_Pos < 10'd328)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd443) && (X_Pos < 10'd482) && (Y_Pos > 10'd324) && (Y_Pos < 10'd328)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd324) && (Y_Pos < 10'd328)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd324) && (Y_Pos < 10'd328)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd325) && (Y_Pos < 10'd329)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd325) && (Y_Pos < 10'd329)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd156) && (X_Pos < 10'd161) && (Y_Pos > 10'd325) && (Y_Pos < 10'd329)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd193) && (X_Pos < 10'd198) && (Y_Pos > 10'd325) && (Y_Pos < 10'd329)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd227) && (X_Pos < 10'd232) && (Y_Pos > 10'd325) && (Y_Pos < 10'd329)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd278) && (X_Pos < 10'd283) && (Y_Pos > 10'd325) && (Y_Pos < 10'd329)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd325) && (Y_Pos < 10'd329)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd325) && (Y_Pos < 10'd329)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd356) && (X_Pos < 10'd361) && (Y_Pos > 10'd325) && (Y_Pos < 10'd329)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd407) && (X_Pos < 10'd412) && (Y_Pos > 10'd325) && (Y_Pos < 10'd329)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd441) && (X_Pos < 10'd446) && (Y_Pos > 10'd325) && (Y_Pos < 10'd329)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd478) && (X_Pos < 10'd483) && (Y_Pos > 10'd325) && (Y_Pos < 10'd329)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd325) && (Y_Pos < 10'd329)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd325) && (Y_Pos < 10'd329)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd326) && (Y_Pos < 10'd330)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd326) && (Y_Pos < 10'd330)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd155) && (X_Pos < 10'd160) && (Y_Pos > 10'd326) && (Y_Pos < 10'd330)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd193) && (X_Pos < 10'd198) && (Y_Pos > 10'd326) && (Y_Pos < 10'd330)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd226) && (X_Pos < 10'd231) && (Y_Pos > 10'd326) && (Y_Pos < 10'd330)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd279) && (X_Pos < 10'd284) && (Y_Pos > 10'd326) && (Y_Pos < 10'd330)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd326) && (Y_Pos < 10'd330)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd326) && (Y_Pos < 10'd330)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd355) && (X_Pos < 10'd360) && (Y_Pos > 10'd326) && (Y_Pos < 10'd330)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd408) && (X_Pos < 10'd413) && (Y_Pos > 10'd326) && (Y_Pos < 10'd330)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd441) && (X_Pos < 10'd446) && (Y_Pos > 10'd326) && (Y_Pos < 10'd330)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd479) && (X_Pos < 10'd484) && (Y_Pos > 10'd326) && (Y_Pos < 10'd330)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd326) && (Y_Pos < 10'd330)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd326) && (Y_Pos < 10'd330)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd327) && (Y_Pos < 10'd331)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd327) && (Y_Pos < 10'd331)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd154) && (X_Pos < 10'd159) && (Y_Pos > 10'd327) && (Y_Pos < 10'd331)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd327) && (Y_Pos < 10'd331)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd327) && (Y_Pos < 10'd331)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd280) && (X_Pos < 10'd285) && (Y_Pos > 10'd327) && (Y_Pos < 10'd331)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd327) && (Y_Pos < 10'd331)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd327) && (Y_Pos < 10'd331)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd354) && (X_Pos < 10'd359) && (Y_Pos > 10'd327) && (Y_Pos < 10'd331)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd327) && (Y_Pos < 10'd331)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd327) && (Y_Pos < 10'd331)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd480) && (X_Pos < 10'd485) && (Y_Pos > 10'd327) && (Y_Pos < 10'd331)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd327) && (Y_Pos < 10'd331)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd327) && (Y_Pos < 10'd331)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd328) && (Y_Pos < 10'd332)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd328) && (Y_Pos < 10'd332)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd154) && (X_Pos < 10'd159) && (Y_Pos > 10'd328) && (Y_Pos < 10'd332)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd328) && (Y_Pos < 10'd332)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd328) && (Y_Pos < 10'd332)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd280) && (X_Pos < 10'd285) && (Y_Pos > 10'd328) && (Y_Pos < 10'd332)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd328) && (Y_Pos < 10'd332)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd328) && (Y_Pos < 10'd332)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd354) && (X_Pos < 10'd359) && (Y_Pos > 10'd328) && (Y_Pos < 10'd332)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd328) && (Y_Pos < 10'd332)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd328) && (Y_Pos < 10'd332)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd480) && (X_Pos < 10'd485) && (Y_Pos > 10'd328) && (Y_Pos < 10'd332)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd328) && (Y_Pos < 10'd332)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd328) && (Y_Pos < 10'd332)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd329) && (Y_Pos < 10'd333)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd329) && (Y_Pos < 10'd333)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd154) && (X_Pos < 10'd159) && (Y_Pos > 10'd329) && (Y_Pos < 10'd333)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd329) && (Y_Pos < 10'd333)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd329) && (Y_Pos < 10'd333)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd280) && (X_Pos < 10'd285) && (Y_Pos > 10'd329) && (Y_Pos < 10'd333)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd329) && (Y_Pos < 10'd333)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd329) && (Y_Pos < 10'd333)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd354) && (X_Pos < 10'd359) && (Y_Pos > 10'd329) && (Y_Pos < 10'd333)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd329) && (Y_Pos < 10'd333)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd329) && (Y_Pos < 10'd333)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd480) && (X_Pos < 10'd485) && (Y_Pos > 10'd329) && (Y_Pos < 10'd333)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd329) && (Y_Pos < 10'd333)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd329) && (Y_Pos < 10'd333)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd330) && (Y_Pos < 10'd334)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd330) && (Y_Pos < 10'd334)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd154) && (X_Pos < 10'd159) && (Y_Pos > 10'd330) && (Y_Pos < 10'd334)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd330) && (Y_Pos < 10'd334)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd330) && (Y_Pos < 10'd334)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd280) && (X_Pos < 10'd285) && (Y_Pos > 10'd330) && (Y_Pos < 10'd334)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd330) && (Y_Pos < 10'd334)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd330) && (Y_Pos < 10'd334)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd354) && (X_Pos < 10'd359) && (Y_Pos > 10'd330) && (Y_Pos < 10'd334)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd330) && (Y_Pos < 10'd334)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd330) && (Y_Pos < 10'd334)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd480) && (X_Pos < 10'd485) && (Y_Pos > 10'd330) && (Y_Pos < 10'd334)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd330) && (Y_Pos < 10'd334)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd330) && (Y_Pos < 10'd334)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd331) && (Y_Pos < 10'd335)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd331) && (Y_Pos < 10'd335)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd154) && (X_Pos < 10'd159) && (Y_Pos > 10'd331) && (Y_Pos < 10'd335)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd331) && (Y_Pos < 10'd335)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd331) && (Y_Pos < 10'd335)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd280) && (X_Pos < 10'd285) && (Y_Pos > 10'd331) && (Y_Pos < 10'd335)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd331) && (Y_Pos < 10'd335)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd331) && (Y_Pos < 10'd335)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd354) && (X_Pos < 10'd359) && (Y_Pos > 10'd331) && (Y_Pos < 10'd335)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd331) && (Y_Pos < 10'd335)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd331) && (Y_Pos < 10'd335)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd480) && (X_Pos < 10'd485) && (Y_Pos > 10'd331) && (Y_Pos < 10'd335)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd331) && (Y_Pos < 10'd335)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd331) && (Y_Pos < 10'd335)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd332) && (Y_Pos < 10'd336)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd332) && (Y_Pos < 10'd336)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd154) && (X_Pos < 10'd159) && (Y_Pos > 10'd332) && (Y_Pos < 10'd336)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd332) && (Y_Pos < 10'd336)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd332) && (Y_Pos < 10'd336)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd280) && (X_Pos < 10'd285) && (Y_Pos > 10'd332) && (Y_Pos < 10'd336)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd332) && (Y_Pos < 10'd336)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd332) && (Y_Pos < 10'd336)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd354) && (X_Pos < 10'd359) && (Y_Pos > 10'd332) && (Y_Pos < 10'd336)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd332) && (Y_Pos < 10'd336)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd332) && (Y_Pos < 10'd336)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd480) && (X_Pos < 10'd485) && (Y_Pos > 10'd332) && (Y_Pos < 10'd336)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd332) && (Y_Pos < 10'd336)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd332) && (Y_Pos < 10'd336)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd333) && (Y_Pos < 10'd337)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd333) && (Y_Pos < 10'd337)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd155) && (X_Pos < 10'd160) && (Y_Pos > 10'd333) && (Y_Pos < 10'd337)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd333) && (Y_Pos < 10'd337)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd227) && (X_Pos < 10'd232) && (Y_Pos > 10'd333) && (Y_Pos < 10'd337)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd279) && (X_Pos < 10'd284) && (Y_Pos > 10'd333) && (Y_Pos < 10'd337)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd312) && (X_Pos < 10'd317) && (Y_Pos > 10'd333) && (Y_Pos < 10'd337)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd322) && (X_Pos < 10'd327) && (Y_Pos > 10'd333) && (Y_Pos < 10'd337)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd355) && (X_Pos < 10'd360) && (Y_Pos > 10'd333) && (Y_Pos < 10'd337)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd407) && (X_Pos < 10'd412) && (Y_Pos > 10'd333) && (Y_Pos < 10'd337)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd333) && (Y_Pos < 10'd337)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd479) && (X_Pos < 10'd484) && (Y_Pos > 10'd333) && (Y_Pos < 10'd337)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd333) && (Y_Pos < 10'd337)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd333) && (Y_Pos < 10'd337)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd334) && (Y_Pos < 10'd338)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd334) && (Y_Pos < 10'd338)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd156) && (X_Pos < 10'd161) && (Y_Pos > 10'd334) && (Y_Pos < 10'd338)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd334) && (Y_Pos < 10'd338)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd227) && (X_Pos < 10'd232) && (Y_Pos > 10'd334) && (Y_Pos < 10'd338)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd278) && (X_Pos < 10'd283) && (Y_Pos > 10'd334) && (Y_Pos < 10'd338)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd313) && (X_Pos < 10'd318) && (Y_Pos > 10'd334) && (Y_Pos < 10'd338)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd321) && (X_Pos < 10'd326) && (Y_Pos > 10'd334) && (Y_Pos < 10'd338)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd356) && (X_Pos < 10'd361) && (Y_Pos > 10'd334) && (Y_Pos < 10'd338)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd407) && (X_Pos < 10'd412) && (Y_Pos > 10'd334) && (Y_Pos < 10'd338)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd334) && (Y_Pos < 10'd338)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd478) && (X_Pos < 10'd483) && (Y_Pos > 10'd334) && (Y_Pos < 10'd338)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd334) && (Y_Pos < 10'd338)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd334) && (Y_Pos < 10'd338)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd335) && (Y_Pos < 10'd339)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd335) && (Y_Pos < 10'd339)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd157) && (X_Pos < 10'd183) && (Y_Pos > 10'd335) && (Y_Pos < 10'd339)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd335) && (Y_Pos < 10'd339)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd229) && (X_Pos < 10'd282) && (Y_Pos > 10'd335) && (Y_Pos < 10'd339)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd314) && (X_Pos < 10'd325) && (Y_Pos > 10'd335) && (Y_Pos < 10'd339)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd357) && (X_Pos < 10'd410) && (Y_Pos > 10'd335) && (Y_Pos < 10'd339)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd335) && (Y_Pos < 10'd339)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd456) && (X_Pos < 10'd482) && (Y_Pos > 10'd335) && (Y_Pos < 10'd339)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd335) && (Y_Pos < 10'd339)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd335) && (Y_Pos < 10'd339)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd336) && (Y_Pos < 10'd340)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd336) && (Y_Pos < 10'd340)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd180) && (X_Pos < 10'd185) && (Y_Pos > 10'd336) && (Y_Pos < 10'd340)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd336) && (Y_Pos < 10'd340)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd336) && (Y_Pos < 10'd340)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd454) && (X_Pos < 10'd459) && (Y_Pos > 10'd336) && (Y_Pos < 10'd340)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd336) && (Y_Pos < 10'd340)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd336) && (Y_Pos < 10'd340)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd337) && (Y_Pos < 10'd341)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd337) && (Y_Pos < 10'd341)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd181) && (X_Pos < 10'd186) && (Y_Pos > 10'd337) && (Y_Pos < 10'd341)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd337) && (Y_Pos < 10'd341)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd337) && (Y_Pos < 10'd341)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd453) && (X_Pos < 10'd458) && (Y_Pos > 10'd337) && (Y_Pos < 10'd341)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd337) && (Y_Pos < 10'd341)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd337) && (Y_Pos < 10'd341)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd338) && (Y_Pos < 10'd342)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd338) && (Y_Pos < 10'd342)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd182) && (X_Pos < 10'd187) && (Y_Pos > 10'd338) && (Y_Pos < 10'd342)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd338) && (Y_Pos < 10'd342)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd338) && (Y_Pos < 10'd342)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd452) && (X_Pos < 10'd457) && (Y_Pos > 10'd338) && (Y_Pos < 10'd342)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd338) && (Y_Pos < 10'd342)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd338) && (Y_Pos < 10'd342)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd339) && (Y_Pos < 10'd343)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd339) && (Y_Pos < 10'd343)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd182) && (X_Pos < 10'd187) && (Y_Pos > 10'd339) && (Y_Pos < 10'd343)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd339) && (Y_Pos < 10'd343)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd339) && (Y_Pos < 10'd343)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd452) && (X_Pos < 10'd457) && (Y_Pos > 10'd339) && (Y_Pos < 10'd343)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd339) && (Y_Pos < 10'd343)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd339) && (Y_Pos < 10'd343)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd340) && (Y_Pos < 10'd344)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd340) && (Y_Pos < 10'd344)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd182) && (X_Pos < 10'd187) && (Y_Pos > 10'd340) && (Y_Pos < 10'd344)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd340) && (Y_Pos < 10'd344)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd340) && (Y_Pos < 10'd344)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd452) && (X_Pos < 10'd457) && (Y_Pos > 10'd340) && (Y_Pos < 10'd344)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd340) && (Y_Pos < 10'd344)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd340) && (Y_Pos < 10'd344)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd341) && (Y_Pos < 10'd345)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd341) && (Y_Pos < 10'd345)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd182) && (X_Pos < 10'd187) && (Y_Pos > 10'd341) && (Y_Pos < 10'd345)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd341) && (Y_Pos < 10'd345)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd341) && (Y_Pos < 10'd345)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd452) && (X_Pos < 10'd457) && (Y_Pos > 10'd341) && (Y_Pos < 10'd345)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd341) && (Y_Pos < 10'd345)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd341) && (Y_Pos < 10'd345)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd342) && (Y_Pos < 10'd346)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd342) && (Y_Pos < 10'd346)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd182) && (X_Pos < 10'd187) && (Y_Pos > 10'd342) && (Y_Pos < 10'd346)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd342) && (Y_Pos < 10'd346)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd342) && (Y_Pos < 10'd346)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd452) && (X_Pos < 10'd457) && (Y_Pos > 10'd342) && (Y_Pos < 10'd346)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd342) && (Y_Pos < 10'd346)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd342) && (Y_Pos < 10'd346)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd343) && (Y_Pos < 10'd347)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd343) && (Y_Pos < 10'd347)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd182) && (X_Pos < 10'd187) && (Y_Pos > 10'd343) && (Y_Pos < 10'd347)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd343) && (Y_Pos < 10'd347)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd343) && (Y_Pos < 10'd347)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd452) && (X_Pos < 10'd457) && (Y_Pos > 10'd343) && (Y_Pos < 10'd347)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd343) && (Y_Pos < 10'd347)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd343) && (Y_Pos < 10'd347)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd344) && (Y_Pos < 10'd348)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd344) && (Y_Pos < 10'd348)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd182) && (X_Pos < 10'd187) && (Y_Pos > 10'd344) && (Y_Pos < 10'd348)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd344) && (Y_Pos < 10'd348)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd344) && (Y_Pos < 10'd348)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd452) && (X_Pos < 10'd457) && (Y_Pos > 10'd344) && (Y_Pos < 10'd348)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd344) && (Y_Pos < 10'd348)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd344) && (Y_Pos < 10'd348)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd345) && (Y_Pos < 10'd349)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd345) && (Y_Pos < 10'd349)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd182) && (X_Pos < 10'd187) && (Y_Pos > 10'd345) && (Y_Pos < 10'd349)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd345) && (Y_Pos < 10'd349)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd345) && (Y_Pos < 10'd349)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd452) && (X_Pos < 10'd457) && (Y_Pos > 10'd345) && (Y_Pos < 10'd349)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd345) && (Y_Pos < 10'd349)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd345) && (Y_Pos < 10'd349)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd346) && (Y_Pos < 10'd350)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd346) && (Y_Pos < 10'd350)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd182) && (X_Pos < 10'd187) && (Y_Pos > 10'd346) && (Y_Pos < 10'd350)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd346) && (Y_Pos < 10'd350)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd346) && (Y_Pos < 10'd350)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd452) && (X_Pos < 10'd457) && (Y_Pos > 10'd346) && (Y_Pos < 10'd350)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd346) && (Y_Pos < 10'd350)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd346) && (Y_Pos < 10'd350)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd347) && (Y_Pos < 10'd351)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd347) && (Y_Pos < 10'd351)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd182) && (X_Pos < 10'd187) && (Y_Pos > 10'd347) && (Y_Pos < 10'd351)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd347) && (Y_Pos < 10'd351)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd347) && (Y_Pos < 10'd351)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd452) && (X_Pos < 10'd457) && (Y_Pos > 10'd347) && (Y_Pos < 10'd351)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd347) && (Y_Pos < 10'd351)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd347) && (Y_Pos < 10'd351)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd348) && (Y_Pos < 10'd352)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd348) && (Y_Pos < 10'd352)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd182) && (X_Pos < 10'd187) && (Y_Pos > 10'd348) && (Y_Pos < 10'd352)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd348) && (Y_Pos < 10'd352)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd348) && (Y_Pos < 10'd352)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd452) && (X_Pos < 10'd457) && (Y_Pos > 10'd348) && (Y_Pos < 10'd352)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd348) && (Y_Pos < 10'd352)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd348) && (Y_Pos < 10'd352)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd349) && (Y_Pos < 10'd353)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd349) && (Y_Pos < 10'd353)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd182) && (X_Pos < 10'd187) && (Y_Pos > 10'd349) && (Y_Pos < 10'd353)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd349) && (Y_Pos < 10'd353)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd349) && (Y_Pos < 10'd353)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd452) && (X_Pos < 10'd457) && (Y_Pos > 10'd349) && (Y_Pos < 10'd353)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd349) && (Y_Pos < 10'd353)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd349) && (Y_Pos < 10'd353)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd350) && (Y_Pos < 10'd354)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd350) && (Y_Pos < 10'd354)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd182) && (X_Pos < 10'd187) && (Y_Pos > 10'd350) && (Y_Pos < 10'd354)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd350) && (Y_Pos < 10'd354)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd350) && (Y_Pos < 10'd354)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd452) && (X_Pos < 10'd457) && (Y_Pos > 10'd350) && (Y_Pos < 10'd354)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd350) && (Y_Pos < 10'd354)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd350) && (Y_Pos < 10'd354)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd351) && (Y_Pos < 10'd355)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd351) && (Y_Pos < 10'd355)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd182) && (X_Pos < 10'd187) && (Y_Pos > 10'd351) && (Y_Pos < 10'd355)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd351) && (Y_Pos < 10'd355)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd351) && (Y_Pos < 10'd355)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd452) && (X_Pos < 10'd457) && (Y_Pos > 10'd351) && (Y_Pos < 10'd355)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd351) && (Y_Pos < 10'd355)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd351) && (Y_Pos < 10'd355)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd352) && (Y_Pos < 10'd356)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd352) && (Y_Pos < 10'd356)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd182) && (X_Pos < 10'd187) && (Y_Pos > 10'd352) && (Y_Pos < 10'd356)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd352) && (Y_Pos < 10'd356)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd352) && (Y_Pos < 10'd356)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd452) && (X_Pos < 10'd457) && (Y_Pos > 10'd352) && (Y_Pos < 10'd356)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd352) && (Y_Pos < 10'd356)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd352) && (Y_Pos < 10'd356)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd353) && (Y_Pos < 10'd357)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd353) && (Y_Pos < 10'd357)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd182) && (X_Pos < 10'd187) && (Y_Pos > 10'd353) && (Y_Pos < 10'd357)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd353) && (Y_Pos < 10'd357)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd353) && (Y_Pos < 10'd357)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd452) && (X_Pos < 10'd457) && (Y_Pos > 10'd353) && (Y_Pos < 10'd357)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd353) && (Y_Pos < 10'd357)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd353) && (Y_Pos < 10'd357)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd354) && (Y_Pos < 10'd358)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd354) && (Y_Pos < 10'd358)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd182) && (X_Pos < 10'd187) && (Y_Pos > 10'd354) && (Y_Pos < 10'd358)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd354) && (Y_Pos < 10'd358)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd354) && (Y_Pos < 10'd358)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd452) && (X_Pos < 10'd457) && (Y_Pos > 10'd354) && (Y_Pos < 10'd358)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd354) && (Y_Pos < 10'd358)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd354) && (Y_Pos < 10'd358)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd355) && (Y_Pos < 10'd359)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd355) && (Y_Pos < 10'd359)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd182) && (X_Pos < 10'd187) && (Y_Pos > 10'd355) && (Y_Pos < 10'd359)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd355) && (Y_Pos < 10'd359)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd355) && (Y_Pos < 10'd359)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd452) && (X_Pos < 10'd457) && (Y_Pos > 10'd355) && (Y_Pos < 10'd359)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd355) && (Y_Pos < 10'd359)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd355) && (Y_Pos < 10'd359)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd356) && (Y_Pos < 10'd360)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd356) && (Y_Pos < 10'd360)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd182) && (X_Pos < 10'd187) && (Y_Pos > 10'd356) && (Y_Pos < 10'd360)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd356) && (Y_Pos < 10'd360)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd356) && (Y_Pos < 10'd360)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd452) && (X_Pos < 10'd457) && (Y_Pos > 10'd356) && (Y_Pos < 10'd360)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd356) && (Y_Pos < 10'd360)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd356) && (Y_Pos < 10'd360)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd357) && (Y_Pos < 10'd361)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd357) && (Y_Pos < 10'd361)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd182) && (X_Pos < 10'd187) && (Y_Pos > 10'd357) && (Y_Pos < 10'd361)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd357) && (Y_Pos < 10'd361)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd357) && (Y_Pos < 10'd361)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd452) && (X_Pos < 10'd457) && (Y_Pos > 10'd357) && (Y_Pos < 10'd361)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd357) && (Y_Pos < 10'd361)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd357) && (Y_Pos < 10'd361)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd358) && (Y_Pos < 10'd362)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd358) && (Y_Pos < 10'd362)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd182) && (X_Pos < 10'd187) && (Y_Pos > 10'd358) && (Y_Pos < 10'd362)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd358) && (Y_Pos < 10'd362)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd358) && (Y_Pos < 10'd362)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd452) && (X_Pos < 10'd457) && (Y_Pos > 10'd358) && (Y_Pos < 10'd362)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd358) && (Y_Pos < 10'd362)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd358) && (Y_Pos < 10'd362)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd359) && (Y_Pos < 10'd363)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd359) && (Y_Pos < 10'd363)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd182) && (X_Pos < 10'd187) && (Y_Pos > 10'd359) && (Y_Pos < 10'd363)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd359) && (Y_Pos < 10'd363)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd359) && (Y_Pos < 10'd363)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd452) && (X_Pos < 10'd457) && (Y_Pos > 10'd359) && (Y_Pos < 10'd363)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd359) && (Y_Pos < 10'd363)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd359) && (Y_Pos < 10'd363)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd360) && (Y_Pos < 10'd364)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd124) && (X_Pos < 10'd129) && (Y_Pos > 10'd360) && (Y_Pos < 10'd364)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd182) && (X_Pos < 10'd187) && (Y_Pos > 10'd360) && (Y_Pos < 10'd364)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd360) && (Y_Pos < 10'd364)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd360) && (Y_Pos < 10'd364)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd452) && (X_Pos < 10'd457) && (Y_Pos > 10'd360) && (Y_Pos < 10'd364)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd510) && (X_Pos < 10'd515) && (Y_Pos > 10'd360) && (Y_Pos < 10'd364)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd360) && (Y_Pos < 10'd364)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd361) && (Y_Pos < 10'd365)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd125) && (X_Pos < 10'd130) && (Y_Pos > 10'd361) && (Y_Pos < 10'd365)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd182) && (X_Pos < 10'd187) && (Y_Pos > 10'd361) && (Y_Pos < 10'd365)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd361) && (Y_Pos < 10'd365)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd361) && (Y_Pos < 10'd365)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd452) && (X_Pos < 10'd457) && (Y_Pos > 10'd361) && (Y_Pos < 10'd365)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd509) && (X_Pos < 10'd514) && (Y_Pos > 10'd361) && (Y_Pos < 10'd365)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd361) && (Y_Pos < 10'd365)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd362) && (Y_Pos < 10'd366)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd127) && (X_Pos < 10'd153) && (Y_Pos > 10'd362) && (Y_Pos < 10'd366)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd182) && (X_Pos < 10'd187) && (Y_Pos > 10'd362) && (Y_Pos < 10'd366)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd362) && (Y_Pos < 10'd366)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd229) && (X_Pos < 10'd239) && (Y_Pos > 10'd362) && (Y_Pos < 10'd366)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd272) && (X_Pos < 10'd367) && (Y_Pos > 10'd362) && (Y_Pos < 10'd366)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd400) && (X_Pos < 10'd410) && (Y_Pos > 10'd362) && (Y_Pos < 10'd366)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd362) && (Y_Pos < 10'd366)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd452) && (X_Pos < 10'd457) && (Y_Pos > 10'd362) && (Y_Pos < 10'd366)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd486) && (X_Pos < 10'd512) && (Y_Pos > 10'd362) && (Y_Pos < 10'd366)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd362) && (Y_Pos < 10'd366)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd363) && (Y_Pos < 10'd367)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd127) && (X_Pos < 10'd154) && (Y_Pos > 10'd363) && (Y_Pos < 10'd367)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd182) && (X_Pos < 10'd187) && (Y_Pos > 10'd363) && (Y_Pos < 10'd367)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd363) && (Y_Pos < 10'd367)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd228) && (X_Pos < 10'd239) && (Y_Pos > 10'd363) && (Y_Pos < 10'd367)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd271) && (X_Pos < 10'd368) && (Y_Pos > 10'd363) && (Y_Pos < 10'd367)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd400) && (X_Pos < 10'd411) && (Y_Pos > 10'd363) && (Y_Pos < 10'd367)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd363) && (Y_Pos < 10'd367)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd452) && (X_Pos < 10'd457) && (Y_Pos > 10'd363) && (Y_Pos < 10'd367)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd485) && (X_Pos < 10'd512) && (Y_Pos > 10'd363) && (Y_Pos < 10'd367)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd363) && (Y_Pos < 10'd367)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd364) && (Y_Pos < 10'd368)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd150) && (X_Pos < 10'd155) && (Y_Pos > 10'd364) && (Y_Pos < 10'd368)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd182) && (X_Pos < 10'd187) && (Y_Pos > 10'd364) && (Y_Pos < 10'd368)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd364) && (Y_Pos < 10'd368)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd227) && (X_Pos < 10'd232) && (Y_Pos > 10'd364) && (Y_Pos < 10'd368)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd236) && (X_Pos < 10'd241) && (Y_Pos > 10'd364) && (Y_Pos < 10'd368)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd270) && (X_Pos < 10'd275) && (Y_Pos > 10'd364) && (Y_Pos < 10'd368)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd364) && (X_Pos < 10'd369) && (Y_Pos > 10'd364) && (Y_Pos < 10'd368)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd398) && (X_Pos < 10'd403) && (Y_Pos > 10'd364) && (Y_Pos < 10'd368)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd407) && (X_Pos < 10'd412) && (Y_Pos > 10'd364) && (Y_Pos < 10'd368)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd364) && (Y_Pos < 10'd368)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd452) && (X_Pos < 10'd457) && (Y_Pos > 10'd364) && (Y_Pos < 10'd368)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd484) && (X_Pos < 10'd489) && (Y_Pos > 10'd364) && (Y_Pos < 10'd368)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd364) && (Y_Pos < 10'd368)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd365) && (Y_Pos < 10'd369)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd151) && (X_Pos < 10'd156) && (Y_Pos > 10'd365) && (Y_Pos < 10'd369)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd182) && (X_Pos < 10'd187) && (Y_Pos > 10'd365) && (Y_Pos < 10'd369)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd365) && (Y_Pos < 10'd369)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd231) && (Y_Pos > 10'd365) && (Y_Pos < 10'd369)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd237) && (X_Pos < 10'd242) && (Y_Pos > 10'd365) && (Y_Pos < 10'd369)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd274) && (Y_Pos > 10'd365) && (Y_Pos < 10'd369)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd365) && (X_Pos < 10'd371) && (Y_Pos > 10'd365) && (Y_Pos < 10'd369)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd397) && (X_Pos < 10'd402) && (Y_Pos > 10'd365) && (Y_Pos < 10'd369)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd408) && (X_Pos < 10'd414) && (Y_Pos > 10'd365) && (Y_Pos < 10'd369)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd365) && (Y_Pos < 10'd369)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd452) && (X_Pos < 10'd457) && (Y_Pos > 10'd365) && (Y_Pos < 10'd369)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd483) && (X_Pos < 10'd488) && (Y_Pos > 10'd365) && (Y_Pos < 10'd369)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd365) && (Y_Pos < 10'd369)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd366) && (Y_Pos < 10'd370)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd152) && (X_Pos < 10'd157) && (Y_Pos > 10'd366) && (Y_Pos < 10'd370)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd182) && (X_Pos < 10'd187) && (Y_Pos > 10'd366) && (Y_Pos < 10'd370)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd366) && (Y_Pos < 10'd370)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd366) && (Y_Pos < 10'd370)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd366) && (Y_Pos < 10'd370)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd366) && (Y_Pos < 10'd370)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd366) && (Y_Pos < 10'd370)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd366) && (Y_Pos < 10'd370)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd366) && (Y_Pos < 10'd370)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd366) && (Y_Pos < 10'd370)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd452) && (X_Pos < 10'd457) && (Y_Pos > 10'd366) && (Y_Pos < 10'd370)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd482) && (X_Pos < 10'd487) && (Y_Pos > 10'd366) && (Y_Pos < 10'd370)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd366) && (Y_Pos < 10'd370)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd367) && (Y_Pos < 10'd371)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd152) && (X_Pos < 10'd157) && (Y_Pos > 10'd367) && (Y_Pos < 10'd371)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd182) && (X_Pos < 10'd187) && (Y_Pos > 10'd367) && (Y_Pos < 10'd371)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd367) && (Y_Pos < 10'd371)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd367) && (Y_Pos < 10'd371)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd367) && (Y_Pos < 10'd371)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd367) && (Y_Pos < 10'd371)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd367) && (Y_Pos < 10'd371)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd367) && (Y_Pos < 10'd371)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd367) && (Y_Pos < 10'd371)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd367) && (Y_Pos < 10'd371)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd452) && (X_Pos < 10'd457) && (Y_Pos > 10'd367) && (Y_Pos < 10'd371)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd482) && (X_Pos < 10'd487) && (Y_Pos > 10'd367) && (Y_Pos < 10'd371)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd367) && (Y_Pos < 10'd371)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd368) && (Y_Pos < 10'd372)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd152) && (X_Pos < 10'd157) && (Y_Pos > 10'd368) && (Y_Pos < 10'd372)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd182) && (X_Pos < 10'd187) && (Y_Pos > 10'd368) && (Y_Pos < 10'd372)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd368) && (Y_Pos < 10'd372)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd368) && (Y_Pos < 10'd372)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd368) && (Y_Pos < 10'd372)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd368) && (Y_Pos < 10'd372)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd368) && (Y_Pos < 10'd372)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd368) && (Y_Pos < 10'd372)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd368) && (Y_Pos < 10'd372)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd368) && (Y_Pos < 10'd372)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd452) && (X_Pos < 10'd457) && (Y_Pos > 10'd368) && (Y_Pos < 10'd372)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd482) && (X_Pos < 10'd487) && (Y_Pos > 10'd368) && (Y_Pos < 10'd372)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd368) && (Y_Pos < 10'd372)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd369) && (Y_Pos < 10'd373)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd152) && (X_Pos < 10'd157) && (Y_Pos > 10'd369) && (Y_Pos < 10'd373)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd182) && (X_Pos < 10'd187) && (Y_Pos > 10'd369) && (Y_Pos < 10'd373)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd369) && (Y_Pos < 10'd373)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd369) && (Y_Pos < 10'd373)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd369) && (Y_Pos < 10'd373)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd369) && (Y_Pos < 10'd373)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd369) && (Y_Pos < 10'd373)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd369) && (Y_Pos < 10'd373)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd369) && (Y_Pos < 10'd373)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd369) && (Y_Pos < 10'd373)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd452) && (X_Pos < 10'd457) && (Y_Pos > 10'd369) && (Y_Pos < 10'd373)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd482) && (X_Pos < 10'd487) && (Y_Pos > 10'd369) && (Y_Pos < 10'd373)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd369) && (Y_Pos < 10'd373)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd370) && (Y_Pos < 10'd374)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd152) && (X_Pos < 10'd157) && (Y_Pos > 10'd370) && (Y_Pos < 10'd374)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd182) && (X_Pos < 10'd187) && (Y_Pos > 10'd370) && (Y_Pos < 10'd374)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd370) && (Y_Pos < 10'd374)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd370) && (Y_Pos < 10'd374)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd370) && (Y_Pos < 10'd374)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd370) && (Y_Pos < 10'd374)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd370) && (Y_Pos < 10'd374)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd370) && (Y_Pos < 10'd374)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd370) && (Y_Pos < 10'd374)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd370) && (Y_Pos < 10'd374)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd452) && (X_Pos < 10'd457) && (Y_Pos > 10'd370) && (Y_Pos < 10'd374)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd482) && (X_Pos < 10'd487) && (Y_Pos > 10'd370) && (Y_Pos < 10'd374)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd370) && (Y_Pos < 10'd374)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd371) && (Y_Pos < 10'd375)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd151) && (X_Pos < 10'd157) && (Y_Pos > 10'd371) && (Y_Pos < 10'd375)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd182) && (X_Pos < 10'd188) && (Y_Pos > 10'd371) && (Y_Pos < 10'd375)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd194) && (X_Pos < 10'd199) && (Y_Pos > 10'd371) && (Y_Pos < 10'd375)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd371) && (Y_Pos < 10'd375)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd371) && (Y_Pos < 10'd375)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd371) && (Y_Pos < 10'd375)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd371) && (Y_Pos < 10'd375)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd371) && (Y_Pos < 10'd375)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd371) && (Y_Pos < 10'd375)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd440) && (X_Pos < 10'd445) && (Y_Pos > 10'd371) && (Y_Pos < 10'd375)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd451) && (X_Pos < 10'd457) && (Y_Pos > 10'd371) && (Y_Pos < 10'd375)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd482) && (X_Pos < 10'd488) && (Y_Pos > 10'd371) && (Y_Pos < 10'd375)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd371) && (Y_Pos < 10'd375)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd372) && (Y_Pos < 10'd376)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd150) && (X_Pos < 10'd155) && (Y_Pos > 10'd372) && (Y_Pos < 10'd376)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd184) && (X_Pos < 10'd189) && (Y_Pos > 10'd372) && (Y_Pos < 10'd376)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd193) && (X_Pos < 10'd198) && (Y_Pos > 10'd372) && (Y_Pos < 10'd376)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd372) && (Y_Pos < 10'd376)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd372) && (Y_Pos < 10'd376)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd270) && (X_Pos < 10'd275) && (Y_Pos > 10'd372) && (Y_Pos < 10'd376)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd364) && (X_Pos < 10'd369) && (Y_Pos > 10'd372) && (Y_Pos < 10'd376)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd372) && (Y_Pos < 10'd376)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd372) && (Y_Pos < 10'd376)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd441) && (X_Pos < 10'd446) && (Y_Pos > 10'd372) && (Y_Pos < 10'd376)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd450) && (X_Pos < 10'd455) && (Y_Pos > 10'd372) && (Y_Pos < 10'd376)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd484) && (X_Pos < 10'd489) && (Y_Pos > 10'd372) && (Y_Pos < 10'd376)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd372) && (Y_Pos < 10'd376)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd373) && (Y_Pos < 10'd377)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd127) && (X_Pos < 10'd154) && (Y_Pos > 10'd373) && (Y_Pos < 10'd377)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd185) && (X_Pos < 10'd197) && (Y_Pos > 10'd373) && (Y_Pos < 10'd377)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd373) && (Y_Pos < 10'd377)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd373) && (Y_Pos < 10'd377)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd270) && (X_Pos < 10'd312) && (Y_Pos > 10'd373) && (Y_Pos < 10'd377)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd327) && (X_Pos < 10'd369) && (Y_Pos > 10'd373) && (Y_Pos < 10'd377)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd373) && (Y_Pos < 10'd377)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd373) && (Y_Pos < 10'd377)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd442) && (X_Pos < 10'd454) && (Y_Pos > 10'd373) && (Y_Pos < 10'd377)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd485) && (X_Pos < 10'd512) && (Y_Pos > 10'd373) && (Y_Pos < 10'd377)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd373) && (Y_Pos < 10'd377)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd374) && (Y_Pos < 10'd378)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd127) && (X_Pos < 10'd153) && (Y_Pos > 10'd374) && (Y_Pos < 10'd378)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd186) && (X_Pos < 10'd196) && (Y_Pos > 10'd374) && (Y_Pos < 10'd378)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd374) && (Y_Pos < 10'd378)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd374) && (Y_Pos < 10'd378)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd272) && (X_Pos < 10'd312) && (Y_Pos > 10'd374) && (Y_Pos < 10'd378)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd327) && (X_Pos < 10'd367) && (Y_Pos > 10'd374) && (Y_Pos < 10'd378)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd374) && (Y_Pos < 10'd378)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd374) && (Y_Pos < 10'd378)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd443) && (X_Pos < 10'd453) && (Y_Pos > 10'd374) && (Y_Pos < 10'd378)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd486) && (X_Pos < 10'd512) && (Y_Pos > 10'd374) && (Y_Pos < 10'd378)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd374) && (Y_Pos < 10'd378)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd375) && (Y_Pos < 10'd379)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd125) && (X_Pos < 10'd130) && (Y_Pos > 10'd375) && (Y_Pos < 10'd379)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd375) && (Y_Pos < 10'd379)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd375) && (Y_Pos < 10'd379)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd309) && (X_Pos < 10'd314) && (Y_Pos > 10'd375) && (Y_Pos < 10'd379)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd325) && (X_Pos < 10'd330) && (Y_Pos > 10'd375) && (Y_Pos < 10'd379)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd375) && (Y_Pos < 10'd379)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd375) && (Y_Pos < 10'd379)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd509) && (X_Pos < 10'd514) && (Y_Pos > 10'd375) && (Y_Pos < 10'd379)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd375) && (Y_Pos < 10'd379)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd376) && (Y_Pos < 10'd380)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd125) && (X_Pos < 10'd130) && (Y_Pos > 10'd376) && (Y_Pos < 10'd380)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd376) && (Y_Pos < 10'd380)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd376) && (Y_Pos < 10'd380)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd309) && (X_Pos < 10'd314) && (Y_Pos > 10'd376) && (Y_Pos < 10'd380)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd325) && (X_Pos < 10'd330) && (Y_Pos > 10'd376) && (Y_Pos < 10'd380)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd376) && (Y_Pos < 10'd380)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd376) && (Y_Pos < 10'd380)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd509) && (X_Pos < 10'd514) && (Y_Pos > 10'd376) && (Y_Pos < 10'd380)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd376) && (Y_Pos < 10'd380)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd377) && (Y_Pos < 10'd381)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd377) && (Y_Pos < 10'd381)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd377) && (Y_Pos < 10'd381)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd377) && (Y_Pos < 10'd381)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd377) && (Y_Pos < 10'd381)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd377) && (Y_Pos < 10'd381)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd377) && (Y_Pos < 10'd381)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd377) && (Y_Pos < 10'd381)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd377) && (Y_Pos < 10'd381)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd377) && (Y_Pos < 10'd381)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd378) && (Y_Pos < 10'd382)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd378) && (Y_Pos < 10'd382)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd378) && (Y_Pos < 10'd382)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd378) && (Y_Pos < 10'd382)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd378) && (Y_Pos < 10'd382)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd378) && (Y_Pos < 10'd382)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd378) && (Y_Pos < 10'd382)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd378) && (Y_Pos < 10'd382)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd378) && (Y_Pos < 10'd382)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd378) && (Y_Pos < 10'd382)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd379) && (Y_Pos < 10'd383)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd379) && (Y_Pos < 10'd383)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd379) && (Y_Pos < 10'd383)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd379) && (Y_Pos < 10'd383)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd379) && (Y_Pos < 10'd383)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd379) && (Y_Pos < 10'd383)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd379) && (Y_Pos < 10'd383)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd379) && (Y_Pos < 10'd383)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd379) && (Y_Pos < 10'd383)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd379) && (Y_Pos < 10'd383)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd380) && (Y_Pos < 10'd384)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd380) && (Y_Pos < 10'd384)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd380) && (Y_Pos < 10'd384)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd380) && (Y_Pos < 10'd384)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd380) && (Y_Pos < 10'd384)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd380) && (Y_Pos < 10'd384)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd380) && (Y_Pos < 10'd384)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd380) && (Y_Pos < 10'd384)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd380) && (Y_Pos < 10'd384)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd380) && (Y_Pos < 10'd384)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd381) && (Y_Pos < 10'd385)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd381) && (Y_Pos < 10'd385)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd381) && (Y_Pos < 10'd385)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd381) && (Y_Pos < 10'd385)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd381) && (Y_Pos < 10'd385)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd381) && (Y_Pos < 10'd385)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd381) && (Y_Pos < 10'd385)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd381) && (Y_Pos < 10'd385)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd381) && (Y_Pos < 10'd385)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd381) && (Y_Pos < 10'd385)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd382) && (Y_Pos < 10'd386)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd382) && (Y_Pos < 10'd386)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd382) && (Y_Pos < 10'd386)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd382) && (Y_Pos < 10'd386)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd382) && (Y_Pos < 10'd386)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd382) && (Y_Pos < 10'd386)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd382) && (Y_Pos < 10'd386)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd382) && (Y_Pos < 10'd386)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd382) && (Y_Pos < 10'd386)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd382) && (Y_Pos < 10'd386)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd383) && (Y_Pos < 10'd387)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd383) && (Y_Pos < 10'd387)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd383) && (Y_Pos < 10'd387)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd383) && (Y_Pos < 10'd387)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd383) && (Y_Pos < 10'd387)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd383) && (Y_Pos < 10'd387)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd383) && (Y_Pos < 10'd387)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd383) && (Y_Pos < 10'd387)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd383) && (Y_Pos < 10'd387)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd383) && (Y_Pos < 10'd387)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd384) && (Y_Pos < 10'd388)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd384) && (Y_Pos < 10'd388)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd384) && (Y_Pos < 10'd388)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd384) && (Y_Pos < 10'd388)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd384) && (Y_Pos < 10'd388)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd384) && (Y_Pos < 10'd388)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd384) && (Y_Pos < 10'd388)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd384) && (Y_Pos < 10'd388)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd384) && (Y_Pos < 10'd388)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd384) && (Y_Pos < 10'd388)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd385) && (Y_Pos < 10'd389)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd385) && (Y_Pos < 10'd389)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd385) && (Y_Pos < 10'd389)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd385) && (Y_Pos < 10'd389)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd385) && (Y_Pos < 10'd389)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd385) && (Y_Pos < 10'd389)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd385) && (Y_Pos < 10'd389)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd385) && (Y_Pos < 10'd389)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd385) && (Y_Pos < 10'd389)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd385) && (Y_Pos < 10'd389)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd386) && (Y_Pos < 10'd390)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd386) && (Y_Pos < 10'd390)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd386) && (Y_Pos < 10'd390)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd386) && (Y_Pos < 10'd390)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd386) && (Y_Pos < 10'd390)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd386) && (Y_Pos < 10'd390)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd386) && (Y_Pos < 10'd390)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd386) && (Y_Pos < 10'd390)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd386) && (Y_Pos < 10'd390)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd386) && (Y_Pos < 10'd390)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd387) && (Y_Pos < 10'd391)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd387) && (Y_Pos < 10'd391)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd387) && (Y_Pos < 10'd391)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd387) && (Y_Pos < 10'd391)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd387) && (Y_Pos < 10'd391)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd387) && (Y_Pos < 10'd391)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd387) && (Y_Pos < 10'd391)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd387) && (Y_Pos < 10'd391)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd387) && (Y_Pos < 10'd391)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd387) && (Y_Pos < 10'd391)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd388) && (Y_Pos < 10'd392)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd388) && (Y_Pos < 10'd392)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd388) && (Y_Pos < 10'd392)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd388) && (Y_Pos < 10'd392)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd388) && (Y_Pos < 10'd392)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd388) && (Y_Pos < 10'd392)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd388) && (Y_Pos < 10'd392)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd388) && (Y_Pos < 10'd392)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd388) && (Y_Pos < 10'd392)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd388) && (Y_Pos < 10'd392)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd389) && (Y_Pos < 10'd393)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd389) && (Y_Pos < 10'd393)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd389) && (Y_Pos < 10'd393)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd389) && (Y_Pos < 10'd393)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd389) && (Y_Pos < 10'd393)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd389) && (Y_Pos < 10'd393)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd389) && (Y_Pos < 10'd393)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd389) && (Y_Pos < 10'd393)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd389) && (Y_Pos < 10'd393)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd389) && (Y_Pos < 10'd393)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd390) && (Y_Pos < 10'd394)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd390) && (Y_Pos < 10'd394)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd390) && (Y_Pos < 10'd394)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd390) && (Y_Pos < 10'd394)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd390) && (Y_Pos < 10'd394)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd390) && (Y_Pos < 10'd394)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd390) && (Y_Pos < 10'd394)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd390) && (Y_Pos < 10'd394)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd390) && (Y_Pos < 10'd394)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd390) && (Y_Pos < 10'd394)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd391) && (Y_Pos < 10'd395)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd391) && (Y_Pos < 10'd395)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd391) && (Y_Pos < 10'd395)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd391) && (Y_Pos < 10'd395)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd391) && (Y_Pos < 10'd395)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd391) && (Y_Pos < 10'd395)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd391) && (Y_Pos < 10'd395)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd391) && (Y_Pos < 10'd395)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd391) && (Y_Pos < 10'd395)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd391) && (Y_Pos < 10'd395)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd392) && (Y_Pos < 10'd396)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd392) && (Y_Pos < 10'd396)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd392) && (Y_Pos < 10'd396)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd392) && (Y_Pos < 10'd396)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd392) && (Y_Pos < 10'd396)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd392) && (Y_Pos < 10'd396)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd392) && (Y_Pos < 10'd396)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd392) && (Y_Pos < 10'd396)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd392) && (Y_Pos < 10'd396)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd392) && (Y_Pos < 10'd396)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd393) && (Y_Pos < 10'd397)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd393) && (Y_Pos < 10'd397)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd393) && (Y_Pos < 10'd397)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd393) && (Y_Pos < 10'd397)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd393) && (Y_Pos < 10'd397)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd393) && (Y_Pos < 10'd397)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd393) && (Y_Pos < 10'd397)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd393) && (Y_Pos < 10'd397)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd393) && (Y_Pos < 10'd397)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd393) && (Y_Pos < 10'd397)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd394) && (Y_Pos < 10'd398)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd394) && (Y_Pos < 10'd398)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd394) && (Y_Pos < 10'd398)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd394) && (Y_Pos < 10'd398)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd394) && (Y_Pos < 10'd398)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd394) && (Y_Pos < 10'd398)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd394) && (Y_Pos < 10'd398)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd394) && (Y_Pos < 10'd398)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd394) && (Y_Pos < 10'd398)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd394) && (Y_Pos < 10'd398)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd395) && (Y_Pos < 10'd399)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd395) && (Y_Pos < 10'd399)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd395) && (Y_Pos < 10'd399)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd395) && (Y_Pos < 10'd399)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd395) && (Y_Pos < 10'd399)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd395) && (Y_Pos < 10'd399)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd395) && (Y_Pos < 10'd399)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd395) && (Y_Pos < 10'd399)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd395) && (Y_Pos < 10'd399)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd395) && (Y_Pos < 10'd399)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd396) && (Y_Pos < 10'd400)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd396) && (Y_Pos < 10'd400)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd396) && (Y_Pos < 10'd400)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd396) && (Y_Pos < 10'd400)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd396) && (Y_Pos < 10'd400)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd396) && (Y_Pos < 10'd400)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd396) && (Y_Pos < 10'd400)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd396) && (Y_Pos < 10'd400)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd396) && (Y_Pos < 10'd400)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd396) && (Y_Pos < 10'd400)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd397) && (Y_Pos < 10'd401)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd397) && (Y_Pos < 10'd401)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd397) && (Y_Pos < 10'd401)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd237) && (X_Pos < 10'd243) && (Y_Pos > 10'd397) && (Y_Pos < 10'd401)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd397) && (Y_Pos < 10'd401)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd397) && (Y_Pos < 10'd401)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd402) && (Y_Pos > 10'd397) && (Y_Pos < 10'd401)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd397) && (Y_Pos < 10'd401)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd397) && (Y_Pos < 10'd401)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd397) && (Y_Pos < 10'd401)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd398) && (Y_Pos < 10'd402)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd398) && (Y_Pos < 10'd402)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd398) && (Y_Pos < 10'd402)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd243) && (Y_Pos > 10'd398) && (Y_Pos < 10'd402)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd398) && (Y_Pos < 10'd402)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd398) && (Y_Pos < 10'd402)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd401) && (Y_Pos > 10'd398) && (Y_Pos < 10'd402)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd398) && (Y_Pos < 10'd402)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd398) && (Y_Pos < 10'd402)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd398) && (Y_Pos < 10'd402)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd399) && (Y_Pos < 10'd403)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd399) && (Y_Pos < 10'd403)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd223) && (X_Pos < 10'd229) && (Y_Pos > 10'd399) && (Y_Pos < 10'd403)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd239) && (X_Pos < 10'd244) && (Y_Pos > 10'd399) && (Y_Pos < 10'd403)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd399) && (Y_Pos < 10'd403)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd399) && (Y_Pos < 10'd403)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd395) && (X_Pos < 10'd400) && (Y_Pos > 10'd399) && (Y_Pos < 10'd403)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd410) && (X_Pos < 10'd416) && (Y_Pos > 10'd399) && (Y_Pos < 10'd403)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd399) && (Y_Pos < 10'd403)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd399) && (Y_Pos < 10'd403)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd400) && (Y_Pos < 10'd404)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd400) && (Y_Pos < 10'd404)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd223) && (X_Pos < 10'd228) && (Y_Pos > 10'd400) && (Y_Pos < 10'd404)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd240) && (X_Pos < 10'd245) && (Y_Pos > 10'd400) && (Y_Pos < 10'd404)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd400) && (Y_Pos < 10'd404)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd400) && (Y_Pos < 10'd404)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd394) && (X_Pos < 10'd399) && (Y_Pos > 10'd400) && (Y_Pos < 10'd404)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd411) && (X_Pos < 10'd416) && (Y_Pos > 10'd400) && (Y_Pos < 10'd404)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd400) && (Y_Pos < 10'd404)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd400) && (Y_Pos < 10'd404)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd401) && (Y_Pos < 10'd405)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd401) && (Y_Pos < 10'd405)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd157) && (X_Pos < 10'd226) && (Y_Pos > 10'd401) && (Y_Pos < 10'd405)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd241) && (X_Pos < 10'd282) && (Y_Pos > 10'd401) && (Y_Pos < 10'd405)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd401) && (Y_Pos < 10'd405)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd401) && (Y_Pos < 10'd405)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd357) && (X_Pos < 10'd398) && (Y_Pos > 10'd401) && (Y_Pos < 10'd405)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd413) && (X_Pos < 10'd482) && (Y_Pos > 10'd401) && (Y_Pos < 10'd405)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd401) && (Y_Pos < 10'd405)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd401) && (Y_Pos < 10'd405)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd402) && (Y_Pos < 10'd406)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd402) && (Y_Pos < 10'd406)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd156) && (X_Pos < 10'd226) && (Y_Pos > 10'd402) && (Y_Pos < 10'd406)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd242) && (X_Pos < 10'd283) && (Y_Pos > 10'd402) && (Y_Pos < 10'd406)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd402) && (Y_Pos < 10'd406)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd402) && (Y_Pos < 10'd406)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd356) && (X_Pos < 10'd397) && (Y_Pos > 10'd402) && (Y_Pos < 10'd406)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd413) && (X_Pos < 10'd483) && (Y_Pos > 10'd402) && (Y_Pos < 10'd406)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd402) && (Y_Pos < 10'd406)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd402) && (Y_Pos < 10'd406)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd403) && (Y_Pos < 10'd407)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd403) && (Y_Pos < 10'd407)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd155) && (X_Pos < 10'd160) && (Y_Pos > 10'd403) && (Y_Pos < 10'd407)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd279) && (X_Pos < 10'd284) && (Y_Pos > 10'd403) && (Y_Pos < 10'd407)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd403) && (Y_Pos < 10'd407)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd403) && (Y_Pos < 10'd407)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd355) && (X_Pos < 10'd360) && (Y_Pos > 10'd403) && (Y_Pos < 10'd407)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd479) && (X_Pos < 10'd484) && (Y_Pos > 10'd403) && (Y_Pos < 10'd407)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd403) && (Y_Pos < 10'd407)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd403) && (Y_Pos < 10'd407)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd404) && (Y_Pos < 10'd408)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd404) && (Y_Pos < 10'd408)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd154) && (X_Pos < 10'd159) && (Y_Pos > 10'd404) && (Y_Pos < 10'd408)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd280) && (X_Pos < 10'd285) && (Y_Pos > 10'd404) && (Y_Pos < 10'd408)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd404) && (Y_Pos < 10'd408)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd404) && (Y_Pos < 10'd408)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd354) && (X_Pos < 10'd359) && (Y_Pos > 10'd404) && (Y_Pos < 10'd408)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd480) && (X_Pos < 10'd485) && (Y_Pos > 10'd404) && (Y_Pos < 10'd408)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd404) && (Y_Pos < 10'd408)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd404) && (Y_Pos < 10'd408)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd405) && (Y_Pos < 10'd409)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd405) && (Y_Pos < 10'd409)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd154) && (X_Pos < 10'd159) && (Y_Pos > 10'd405) && (Y_Pos < 10'd409)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd280) && (X_Pos < 10'd285) && (Y_Pos > 10'd405) && (Y_Pos < 10'd409)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd405) && (Y_Pos < 10'd409)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd405) && (Y_Pos < 10'd409)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd354) && (X_Pos < 10'd359) && (Y_Pos > 10'd405) && (Y_Pos < 10'd409)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd480) && (X_Pos < 10'd485) && (Y_Pos > 10'd405) && (Y_Pos < 10'd409)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd405) && (Y_Pos < 10'd409)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd405) && (Y_Pos < 10'd409)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd406) && (Y_Pos < 10'd410)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd406) && (Y_Pos < 10'd410)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd154) && (X_Pos < 10'd159) && (Y_Pos > 10'd406) && (Y_Pos < 10'd410)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd280) && (X_Pos < 10'd285) && (Y_Pos > 10'd406) && (Y_Pos < 10'd410)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd406) && (Y_Pos < 10'd410)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd406) && (Y_Pos < 10'd410)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd354) && (X_Pos < 10'd359) && (Y_Pos > 10'd406) && (Y_Pos < 10'd410)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd480) && (X_Pos < 10'd485) && (Y_Pos > 10'd406) && (Y_Pos < 10'd410)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd406) && (Y_Pos < 10'd410)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd406) && (Y_Pos < 10'd410)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd407) && (Y_Pos < 10'd411)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd407) && (Y_Pos < 10'd411)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd154) && (X_Pos < 10'd159) && (Y_Pos > 10'd407) && (Y_Pos < 10'd411)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd280) && (X_Pos < 10'd285) && (Y_Pos > 10'd407) && (Y_Pos < 10'd411)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd407) && (Y_Pos < 10'd411)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd407) && (Y_Pos < 10'd411)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd354) && (X_Pos < 10'd359) && (Y_Pos > 10'd407) && (Y_Pos < 10'd411)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd480) && (X_Pos < 10'd485) && (Y_Pos > 10'd407) && (Y_Pos < 10'd411)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd407) && (Y_Pos < 10'd411)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd407) && (Y_Pos < 10'd411)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd408) && (Y_Pos < 10'd412)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd408) && (Y_Pos < 10'd412)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd154) && (X_Pos < 10'd159) && (Y_Pos > 10'd408) && (Y_Pos < 10'd412)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd280) && (X_Pos < 10'd285) && (Y_Pos > 10'd408) && (Y_Pos < 10'd412)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd408) && (Y_Pos < 10'd412)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd408) && (Y_Pos < 10'd412)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd354) && (X_Pos < 10'd359) && (Y_Pos > 10'd408) && (Y_Pos < 10'd412)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd480) && (X_Pos < 10'd485) && (Y_Pos > 10'd408) && (Y_Pos < 10'd412)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd408) && (Y_Pos < 10'd412)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd408) && (Y_Pos < 10'd412)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd409) && (Y_Pos < 10'd413)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd409) && (Y_Pos < 10'd413)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd154) && (X_Pos < 10'd159) && (Y_Pos > 10'd409) && (Y_Pos < 10'd413)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd280) && (X_Pos < 10'd285) && (Y_Pos > 10'd409) && (Y_Pos < 10'd413)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd316) && (Y_Pos > 10'd409) && (Y_Pos < 10'd413)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd328) && (Y_Pos > 10'd409) && (Y_Pos < 10'd413)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd354) && (X_Pos < 10'd359) && (Y_Pos > 10'd409) && (Y_Pos < 10'd413)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd480) && (X_Pos < 10'd485) && (Y_Pos > 10'd409) && (Y_Pos < 10'd413)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd409) && (Y_Pos < 10'd413)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd409) && (Y_Pos < 10'd413)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd410) && (Y_Pos < 10'd414)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd410) && (Y_Pos < 10'd414)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd155) && (X_Pos < 10'd160) && (Y_Pos > 10'd410) && (Y_Pos < 10'd414)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd279) && (X_Pos < 10'd284) && (Y_Pos > 10'd410) && (Y_Pos < 10'd414)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd312) && (X_Pos < 10'd317) && (Y_Pos > 10'd410) && (Y_Pos < 10'd414)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd322) && (X_Pos < 10'd327) && (Y_Pos > 10'd410) && (Y_Pos < 10'd414)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd355) && (X_Pos < 10'd360) && (Y_Pos > 10'd410) && (Y_Pos < 10'd414)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd479) && (X_Pos < 10'd484) && (Y_Pos > 10'd410) && (Y_Pos < 10'd414)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd410) && (Y_Pos < 10'd414)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd410) && (Y_Pos < 10'd414)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd411) && (Y_Pos < 10'd415)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd411) && (Y_Pos < 10'd415)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd155) && (X_Pos < 10'd160) && (Y_Pos > 10'd411) && (Y_Pos < 10'd415)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd279) && (X_Pos < 10'd284) && (Y_Pos > 10'd411) && (Y_Pos < 10'd415)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd313) && (X_Pos < 10'd318) && (Y_Pos > 10'd411) && (Y_Pos < 10'd415)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd321) && (X_Pos < 10'd326) && (Y_Pos > 10'd411) && (Y_Pos < 10'd415)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd355) && (X_Pos < 10'd360) && (Y_Pos > 10'd411) && (Y_Pos < 10'd415)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd479) && (X_Pos < 10'd484) && (Y_Pos > 10'd411) && (Y_Pos < 10'd415)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd411) && (Y_Pos < 10'd415)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd411) && (Y_Pos < 10'd415)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd412) && (Y_Pos < 10'd416)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd412) && (Y_Pos < 10'd416)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd157) && (X_Pos < 10'd282) && (Y_Pos > 10'd412) && (Y_Pos < 10'd416)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd314) && (X_Pos < 10'd325) && (Y_Pos > 10'd412) && (Y_Pos < 10'd416)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd357) && (X_Pos < 10'd482) && (Y_Pos > 10'd412) && (Y_Pos < 10'd416)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd412) && (Y_Pos < 10'd416)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd412) && (Y_Pos < 10'd416)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd413) && (Y_Pos < 10'd417)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd413) && (Y_Pos < 10'd417)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd158) && (X_Pos < 10'd281) && (Y_Pos > 10'd413) && (Y_Pos < 10'd417)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd315) && (X_Pos < 10'd324) && (Y_Pos > 10'd413) && (Y_Pos < 10'd417)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd358) && (X_Pos < 10'd481) && (Y_Pos > 10'd413) && (Y_Pos < 10'd417)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd413) && (Y_Pos < 10'd417)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd413) && (Y_Pos < 10'd417)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd414) && (Y_Pos < 10'd418)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd414) && (Y_Pos < 10'd418)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd414) && (Y_Pos < 10'd418)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd414) && (Y_Pos < 10'd418)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd415) && (Y_Pos < 10'd419)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd415) && (Y_Pos < 10'd419)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd415) && (Y_Pos < 10'd419)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd415) && (Y_Pos < 10'd419)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd416) && (Y_Pos < 10'd420)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd416) && (Y_Pos < 10'd420)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd416) && (Y_Pos < 10'd420)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd416) && (Y_Pos < 10'd420)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd417) && (Y_Pos < 10'd421)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd417) && (Y_Pos < 10'd421)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd417) && (Y_Pos < 10'd421)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd417) && (Y_Pos < 10'd421)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd418) && (Y_Pos < 10'd422)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd418) && (Y_Pos < 10'd422)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd418) && (Y_Pos < 10'd422)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd418) && (Y_Pos < 10'd422)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd419) && (Y_Pos < 10'd423)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd419) && (Y_Pos < 10'd423)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd419) && (Y_Pos < 10'd423)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd419) && (Y_Pos < 10'd423)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd420) && (Y_Pos < 10'd424)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd420) && (Y_Pos < 10'd424)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd420) && (Y_Pos < 10'd424)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd420) && (Y_Pos < 10'd424)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd421) && (Y_Pos < 10'd425)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd421) && (Y_Pos < 10'd425)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd421) && (Y_Pos < 10'd425)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd421) && (Y_Pos < 10'd425)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd422) && (Y_Pos < 10'd426)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd422) && (Y_Pos < 10'd426)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd422) && (Y_Pos < 10'd426)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd422) && (Y_Pos < 10'd426)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd423) && (Y_Pos < 10'd427)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd423) && (Y_Pos < 10'd427)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd423) && (Y_Pos < 10'd427)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd423) && (Y_Pos < 10'd427)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd424) && (Y_Pos < 10'd428)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd424) && (Y_Pos < 10'd428)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd424) && (Y_Pos < 10'd428)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd424) && (Y_Pos < 10'd428)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd425) && (Y_Pos < 10'd429)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd425) && (Y_Pos < 10'd429)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd425) && (Y_Pos < 10'd429)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd425) && (Y_Pos < 10'd429)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd426) && (Y_Pos < 10'd430)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd426) && (Y_Pos < 10'd430)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd426) && (Y_Pos < 10'd430)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd426) && (Y_Pos < 10'd430)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd427) && (Y_Pos < 10'd431)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd427) && (Y_Pos < 10'd431)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd427) && (Y_Pos < 10'd431)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd427) && (Y_Pos < 10'd431)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd428) && (Y_Pos < 10'd432)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd428) && (Y_Pos < 10'd432)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd428) && (Y_Pos < 10'd432)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd428) && (Y_Pos < 10'd432)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd429) && (Y_Pos < 10'd433)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd429) && (Y_Pos < 10'd433)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd429) && (Y_Pos < 10'd433)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd429) && (Y_Pos < 10'd433)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd430) && (Y_Pos < 10'd434)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd430) && (Y_Pos < 10'd434)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd430) && (Y_Pos < 10'd434)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd430) && (Y_Pos < 10'd434)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd431) && (Y_Pos < 10'd435)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd431) && (Y_Pos < 10'd435)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd431) && (Y_Pos < 10'd435)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd431) && (Y_Pos < 10'd435)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd432) && (Y_Pos < 10'd436)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd432) && (Y_Pos < 10'd436)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd432) && (Y_Pos < 10'd436)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd432) && (Y_Pos < 10'd436)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd433) && (Y_Pos < 10'd437)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd433) && (Y_Pos < 10'd437)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd433) && (Y_Pos < 10'd437)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd433) && (Y_Pos < 10'd437)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd434) && (Y_Pos < 10'd438)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd434) && (Y_Pos < 10'd438)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd434) && (Y_Pos < 10'd438)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd434) && (Y_Pos < 10'd438)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd435) && (Y_Pos < 10'd439)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd435) && (Y_Pos < 10'd439)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd435) && (Y_Pos < 10'd439)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd435) && (Y_Pos < 10'd439)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd436) && (Y_Pos < 10'd440)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd436) && (Y_Pos < 10'd440)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd436) && (Y_Pos < 10'd440)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd436) && (Y_Pos < 10'd440)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd437) && (Y_Pos < 10'd441)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd437) && (Y_Pos < 10'd441)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd437) && (Y_Pos < 10'd441)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd437) && (Y_Pos < 10'd441)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd438) && (Y_Pos < 10'd442)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd125) && (X_Pos < 10'd130) && (Y_Pos > 10'd438) && (Y_Pos < 10'd442)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd509) && (X_Pos < 10'd514) && (Y_Pos > 10'd438) && (Y_Pos < 10'd442)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd438) && (Y_Pos < 10'd442)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd439) && (Y_Pos < 10'd443)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd125) && (X_Pos < 10'd514) && (Y_Pos > 10'd439) && (Y_Pos < 10'd443)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd439) && (Y_Pos < 10'd443)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd120) && (X_Pos < 10'd125) && (Y_Pos > 10'd440) && (Y_Pos < 10'd444)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd127) && (X_Pos < 10'd512) && (Y_Pos > 10'd440) && (Y_Pos < 10'd444)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd514) && (X_Pos < 10'd519) && (Y_Pos > 10'd440) && (Y_Pos < 10'd444)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd120) && (X_Pos < 10'd125) && (Y_Pos > 10'd441) && (Y_Pos < 10'd445)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd514) && (X_Pos < 10'd519) && (Y_Pos > 10'd441) && (Y_Pos < 10'd445)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd120) && (X_Pos < 10'd125) && (Y_Pos > 10'd442) && (Y_Pos < 10'd446)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd514) && (X_Pos < 10'd519) && (Y_Pos > 10'd442) && (Y_Pos < 10'd446)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd122) && (X_Pos < 10'd128) && (Y_Pos > 10'd443) && (Y_Pos < 10'd447)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd517) && (Y_Pos > 10'd443) && (Y_Pos < 10'd447)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd125) && (X_Pos < 10'd514) && (Y_Pos > 10'd444) && (Y_Pos < 10'd448)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd125) && (X_Pos < 10'd514) && (Y_Pos > 10'd445) && (Y_Pos < 10'd449)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd125) && (X_Pos < 10'd514) && (Y_Pos > 10'd46) && (Y_Pos < 10'd51)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd122) && (X_Pos < 10'd128) && (Y_Pos > 10'd48) && (Y_Pos < 10'd52)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd517) && (Y_Pos > 10'd48) && (Y_Pos < 10'd52)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd120) && (X_Pos < 10'd125) && (Y_Pos > 10'd49) && (Y_Pos < 10'd55)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd514) && (X_Pos < 10'd519) && (Y_Pos > 10'd49) && (Y_Pos < 10'd55)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd127) && (X_Pos < 10'd312) && (Y_Pos > 10'd51) && (Y_Pos < 10'd56)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd327) && (X_Pos < 10'd512) && (Y_Pos > 10'd51) && (Y_Pos < 10'd56)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd125) && (X_Pos < 10'd130) && (Y_Pos > 10'd52) && (Y_Pos < 10'd57)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd309) && (X_Pos < 10'd314) && (Y_Pos > 10'd52) && (Y_Pos < 10'd57)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd325) && (X_Pos < 10'd330) && (Y_Pos > 10'd52) && (Y_Pos < 10'd57)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd509) && (X_Pos < 10'd514) && (Y_Pos > 10'd52) && (Y_Pos < 10'd57)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd52) && (Y_Pos < 10'd172)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd52) && (Y_Pos < 10'd172)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd315) && (Y_Pos > 10'd54) && (Y_Pos < 10'd104)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd324) && (X_Pos < 10'd328) && (Y_Pos > 10'd54) && (Y_Pos < 10'd104)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd312) && (X_Pos < 10'd316) && (Y_Pos > 10'd54) && (Y_Pos < 10'd105)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd327) && (Y_Pos > 10'd54) && (Y_Pos < 10'd105)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd54) && (Y_Pos < 10'd170)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd54) && (Y_Pos < 10'd170)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd158) && (X_Pos < 10'd196) && (Y_Pos > 10'd78) && (Y_Pos < 10'd83)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd229) && (X_Pos < 10'd281) && (Y_Pos > 10'd78) && (Y_Pos < 10'd83)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd358) && (X_Pos < 10'd410) && (Y_Pos > 10'd78) && (Y_Pos < 10'd83)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd443) && (X_Pos < 10'd481) && (Y_Pos > 10'd78) && (Y_Pos < 10'd83)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd228) && (X_Pos < 10'd232) && (Y_Pos > 10'd79) && (Y_Pos < 10'd84)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd407) && (X_Pos < 10'd411) && (Y_Pos > 10'd79) && (Y_Pos < 10'd84)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd157) && (X_Pos < 10'd161) && (Y_Pos > 10'd79) && (Y_Pos < 10'd83)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd278) && (X_Pos < 10'd282) && (Y_Pos > 10'd79) && (Y_Pos < 10'd83)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd357) && (X_Pos < 10'd361) && (Y_Pos > 10'd79) && (Y_Pos < 10'd83)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd478) && (X_Pos < 10'd482) && (Y_Pos > 10'd79) && (Y_Pos < 10'd83)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd156) && (X_Pos < 10'd160) && (Y_Pos > 10'd80) && (Y_Pos < 10'd85)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd193) && (X_Pos < 10'd198) && (Y_Pos > 10'd80) && (Y_Pos < 10'd85)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd227) && (X_Pos < 10'd231) && (Y_Pos > 10'd80) && (Y_Pos < 10'd85)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd279) && (X_Pos < 10'd283) && (Y_Pos > 10'd80) && (Y_Pos < 10'd85)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd356) && (X_Pos < 10'd360) && (Y_Pos > 10'd80) && (Y_Pos < 10'd85)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd408) && (X_Pos < 10'd412) && (Y_Pos > 10'd80) && (Y_Pos < 10'd85)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd441) && (X_Pos < 10'd446) && (Y_Pos > 10'd80) && (Y_Pos < 10'd85)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd479) && (X_Pos < 10'd483) && (Y_Pos > 10'd80) && (Y_Pos < 10'd85)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd155) && (X_Pos < 10'd159) && (Y_Pos > 10'd80) && (Y_Pos < 10'd105)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd280) && (X_Pos < 10'd284) && (Y_Pos > 10'd80) && (Y_Pos < 10'd105)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd355) && (X_Pos < 10'd359) && (Y_Pos > 10'd80) && (Y_Pos < 10'd105)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd480) && (X_Pos < 10'd484) && (Y_Pos > 10'd80) && (Y_Pos < 10'd105)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd199) && (Y_Pos > 10'd81) && (Y_Pos < 10'd104)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd226) && (X_Pos < 10'd230) && (Y_Pos > 10'd81) && (Y_Pos < 10'd104)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd413) && (Y_Pos > 10'd81) && (Y_Pos < 10'd104)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd440) && (X_Pos < 10'd444) && (Y_Pos > 10'd81) && (Y_Pos < 10'd104)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd196) && (X_Pos < 10'd200) && (Y_Pos > 10'd82) && (Y_Pos < 10'd103)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd443) && (Y_Pos > 10'd82) && (Y_Pos < 10'd103)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd154) && (X_Pos < 10'd158) && (Y_Pos > 10'd82) && (Y_Pos < 10'd104)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd229) && (Y_Pos > 10'd82) && (Y_Pos < 10'd104)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd281) && (X_Pos < 10'd285) && (Y_Pos > 10'd82) && (Y_Pos < 10'd104)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd354) && (X_Pos < 10'd358) && (Y_Pos > 10'd82) && (Y_Pos < 10'd104)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd410) && (X_Pos < 10'd414) && (Y_Pos > 10'd82) && (Y_Pos < 10'd104)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd481) && (X_Pos < 10'd485) && (Y_Pos > 10'd82) && (Y_Pos < 10'd104)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd194) && (X_Pos < 10'd198) && (Y_Pos > 10'd100) && (Y_Pos < 10'd105)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd441) && (X_Pos < 10'd445) && (Y_Pos > 10'd100) && (Y_Pos < 10'd105)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd156) && (X_Pos < 10'd160) && (Y_Pos > 10'd101) && (Y_Pos < 10'd106)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd193) && (X_Pos < 10'd197) && (Y_Pos > 10'd101) && (Y_Pos < 10'd106)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd227) && (X_Pos < 10'd232) && (Y_Pos > 10'd101) && (Y_Pos < 10'd106)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd279) && (X_Pos < 10'd283) && (Y_Pos > 10'd101) && (Y_Pos < 10'd106)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd313) && (X_Pos < 10'd318) && (Y_Pos > 10'd101) && (Y_Pos < 10'd106)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd321) && (X_Pos < 10'd326) && (Y_Pos > 10'd101) && (Y_Pos < 10'd106)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd356) && (X_Pos < 10'd360) && (Y_Pos > 10'd101) && (Y_Pos < 10'd106)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd407) && (X_Pos < 10'd412) && (Y_Pos > 10'd101) && (Y_Pos < 10'd106)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd442) && (X_Pos < 10'd446) && (Y_Pos > 10'd101) && (Y_Pos < 10'd106)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd479) && (X_Pos < 10'd483) && (Y_Pos > 10'd101) && (Y_Pos < 10'd106)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd157) && (X_Pos < 10'd196) && (Y_Pos > 10'd102) && (Y_Pos < 10'd107)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd229) && (X_Pos < 10'd282) && (Y_Pos > 10'd102) && (Y_Pos < 10'd107)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd315) && (X_Pos < 10'd324) && (Y_Pos > 10'd102) && (Y_Pos < 10'd107)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd357) && (X_Pos < 10'd410) && (Y_Pos > 10'd102) && (Y_Pos < 10'd107)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd443) && (X_Pos < 10'd482) && (Y_Pos > 10'd102) && (Y_Pos < 10'd107)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd157) && (X_Pos < 10'd196) && (Y_Pos > 10'd130) && (Y_Pos < 10'd135)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd229) && (X_Pos < 10'd239) && (Y_Pos > 10'd130) && (Y_Pos < 10'd135)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd272) && (X_Pos < 10'd367) && (Y_Pos > 10'd130) && (Y_Pos < 10'd135)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd400) && (X_Pos < 10'd410) && (Y_Pos > 10'd130) && (Y_Pos < 10'd135)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd443) && (X_Pos < 10'd482) && (Y_Pos > 10'd130) && (Y_Pos < 10'd135)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd156) && (X_Pos < 10'd160) && (Y_Pos > 10'd131) && (Y_Pos < 10'd136)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd193) && (X_Pos < 10'd197) && (Y_Pos > 10'd131) && (Y_Pos < 10'd136)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd227) && (X_Pos < 10'd232) && (Y_Pos > 10'd131) && (Y_Pos < 10'd136)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd236) && (X_Pos < 10'd240) && (Y_Pos > 10'd131) && (Y_Pos < 10'd136)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd270) && (X_Pos < 10'd275) && (Y_Pos > 10'd131) && (Y_Pos < 10'd136)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd364) && (X_Pos < 10'd369) && (Y_Pos > 10'd131) && (Y_Pos < 10'd136)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd399) && (X_Pos < 10'd403) && (Y_Pos > 10'd131) && (Y_Pos < 10'd136)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd407) && (X_Pos < 10'd412) && (Y_Pos > 10'd131) && (Y_Pos < 10'd136)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd442) && (X_Pos < 10'd446) && (Y_Pos > 10'd131) && (Y_Pos < 10'd136)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd479) && (X_Pos < 10'd483) && (Y_Pos > 10'd131) && (Y_Pos < 10'd136)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd194) && (X_Pos < 10'd198) && (Y_Pos > 10'd132) && (Y_Pos < 10'd137)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd237) && (X_Pos < 10'd241) && (Y_Pos > 10'd132) && (Y_Pos < 10'd137)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd398) && (X_Pos < 10'd402) && (Y_Pos > 10'd132) && (Y_Pos < 10'd137)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd441) && (X_Pos < 10'd445) && (Y_Pos > 10'd132) && (Y_Pos < 10'd137)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd155) && (X_Pos < 10'd159) && (Y_Pos > 10'd132) && (Y_Pos < 10'd144)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd480) && (X_Pos < 10'd484) && (Y_Pos > 10'd132) && (Y_Pos < 10'd144)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd196) && (X_Pos < 10'd200) && (Y_Pos > 10'd133) && (Y_Pos < 10'd142)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd272) && (Y_Pos > 10'd133) && (Y_Pos < 10'd142)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd367) && (X_Pos < 10'd371) && (Y_Pos > 10'd133) && (Y_Pos < 10'd142)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd443) && (Y_Pos > 10'd133) && (Y_Pos < 10'd142)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd154) && (X_Pos < 10'd158) && (Y_Pos > 10'd133) && (Y_Pos < 10'd143)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd199) && (Y_Pos > 10'd133) && (Y_Pos < 10'd143)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd269) && (X_Pos < 10'd273) && (Y_Pos > 10'd133) && (Y_Pos < 10'd143)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd370) && (Y_Pos > 10'd133) && (Y_Pos < 10'd143)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd440) && (X_Pos < 10'd444) && (Y_Pos > 10'd133) && (Y_Pos < 10'd143)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd481) && (X_Pos < 10'd485) && (Y_Pos > 10'd133) && (Y_Pos < 10'd143)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd242) && (Y_Pos > 10'd133) && (Y_Pos < 10'd170)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd397) && (X_Pos < 10'd401) && (Y_Pos > 10'd133) && (Y_Pos < 10'd170)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd230) && (Y_Pos > 10'd133) && (Y_Pos < 10'd220)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd414) && (Y_Pos > 10'd133) && (Y_Pos < 10'd220)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd239) && (X_Pos < 10'd243) && (Y_Pos > 10'd134) && (Y_Pos < 10'd171)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd400) && (Y_Pos > 10'd134) && (Y_Pos < 10'd171)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd156) && (X_Pos < 10'd160) && (Y_Pos > 10'd139) && (Y_Pos < 10'd144)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd194) && (X_Pos < 10'd198) && (Y_Pos > 10'd139) && (Y_Pos < 10'd144)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd270) && (X_Pos < 10'd274) && (Y_Pos > 10'd139) && (Y_Pos < 10'd144)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd365) && (X_Pos < 10'd369) && (Y_Pos > 10'd139) && (Y_Pos < 10'd144)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd441) && (X_Pos < 10'd445) && (Y_Pos > 10'd139) && (Y_Pos < 10'd144)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd479) && (X_Pos < 10'd483) && (Y_Pos > 10'd139) && (Y_Pos < 10'd144)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd193) && (X_Pos < 10'd197) && (Y_Pos > 10'd140) && (Y_Pos < 10'd144)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd442) && (X_Pos < 10'd446) && (Y_Pos > 10'd140) && (Y_Pos < 10'd144)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd271) && (X_Pos < 10'd275) && (Y_Pos > 10'd140) && (Y_Pos < 10'd145)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd364) && (X_Pos < 10'd368) && (Y_Pos > 10'd140) && (Y_Pos < 10'd145)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd157) && (X_Pos < 10'd161) && (Y_Pos > 10'd141) && (Y_Pos < 10'd145)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd478) && (X_Pos < 10'd482) && (Y_Pos > 10'd141) && (Y_Pos < 10'd145)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd158) && (X_Pos < 10'd196) && (Y_Pos > 10'd141) && (Y_Pos < 10'd146)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd272) && (X_Pos < 10'd312) && (Y_Pos > 10'd141) && (Y_Pos < 10'd146)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd327) && (X_Pos < 10'd367) && (Y_Pos > 10'd141) && (Y_Pos < 10'd146)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd443) && (X_Pos < 10'd481) && (Y_Pos > 10'd141) && (Y_Pos < 10'd146)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd309) && (X_Pos < 10'd313) && (Y_Pos > 10'd142) && (Y_Pos < 10'd147)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd326) && (X_Pos < 10'd330) && (Y_Pos > 10'd142) && (Y_Pos < 10'd147)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd310) && (X_Pos < 10'd314) && (Y_Pos > 10'd143) && (Y_Pos < 10'd148)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd325) && (X_Pos < 10'd329) && (Y_Pos > 10'd143) && (Y_Pos < 10'd148)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd315) && (Y_Pos > 10'd144) && (Y_Pos < 10'd181)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd324) && (X_Pos < 10'd328) && (Y_Pos > 10'd144) && (Y_Pos < 10'd181)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd312) && (X_Pos < 10'd316) && (Y_Pos > 10'd145) && (Y_Pos < 10'd182)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd327) && (Y_Pos > 10'd145) && (Y_Pos < 10'd182)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd237) && (X_Pos < 10'd241) && (Y_Pos > 10'd165) && (Y_Pos < 10'd169)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd398) && (X_Pos < 10'd402) && (Y_Pos > 10'd165) && (Y_Pos < 10'd169)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd125) && (X_Pos < 10'd130) && (Y_Pos > 10'd167) && (Y_Pos < 10'd172)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd240) && (X_Pos < 10'd244) && (Y_Pos > 10'd167) && (Y_Pos < 10'd172)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd395) && (X_Pos < 10'd399) && (Y_Pos > 10'd167) && (Y_Pos < 10'd172)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd509) && (X_Pos < 10'd514) && (Y_Pos > 10'd167) && (Y_Pos < 10'd172)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd127) && (X_Pos < 10'd195) && (Y_Pos > 10'd168) && (Y_Pos < 10'd173)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd241) && (X_Pos < 10'd281) && (Y_Pos > 10'd168) && (Y_Pos < 10'd173)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd358) && (X_Pos < 10'd398) && (Y_Pos > 10'd168) && (Y_Pos < 10'd173)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd444) && (X_Pos < 10'd512) && (Y_Pos > 10'd168) && (Y_Pos < 10'd173)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd192) && (X_Pos < 10'd196) && (Y_Pos > 10'd169) && (Y_Pos < 10'd173)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd443) && (X_Pos < 10'd447) && (Y_Pos > 10'd169) && (Y_Pos < 10'd173)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd278) && (X_Pos < 10'd282) && (Y_Pos > 10'd169) && (Y_Pos < 10'd174)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd357) && (X_Pos < 10'd361) && (Y_Pos > 10'd169) && (Y_Pos < 10'd174)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd120) && (X_Pos < 10'd125) && (Y_Pos > 10'd169) && (Y_Pos < 10'd175)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd514) && (X_Pos < 10'd519) && (Y_Pos > 10'd169) && (Y_Pos < 10'd175)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd193) && (X_Pos < 10'd198) && (Y_Pos > 10'd170) && (Y_Pos < 10'd175)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd279) && (X_Pos < 10'd283) && (Y_Pos > 10'd170) && (Y_Pos < 10'd175)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd356) && (X_Pos < 10'd360) && (Y_Pos > 10'd170) && (Y_Pos < 10'd175)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd441) && (X_Pos < 10'd446) && (Y_Pos > 10'd170) && (Y_Pos < 10'd175)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd280) && (X_Pos < 10'd284) && (Y_Pos > 10'd171) && (Y_Pos < 10'd182)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd355) && (X_Pos < 10'd359) && (Y_Pos > 10'd171) && (Y_Pos < 10'd182)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd122) && (X_Pos < 10'd128) && (Y_Pos > 10'd172) && (Y_Pos < 10'd177)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd517) && (Y_Pos > 10'd172) && (Y_Pos < 10'd177)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd281) && (X_Pos < 10'd285) && (Y_Pos > 10'd172) && (Y_Pos < 10'd181)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd354) && (X_Pos < 10'd358) && (Y_Pos > 10'd172) && (Y_Pos < 10'd181)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd200) && (Y_Pos > 10'd172) && (Y_Pos < 10'd220)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd444) && (Y_Pos > 10'd172) && (Y_Pos < 10'd220)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd125) && (X_Pos < 10'd192) && (Y_Pos > 10'd173) && (Y_Pos < 10'd178)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd447) && (X_Pos < 10'd514) && (Y_Pos > 10'd173) && (Y_Pos < 10'd178)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd193) && (Y_Pos > 10'd174) && (Y_Pos < 10'd217)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd446) && (X_Pos < 10'd450) && (Y_Pos > 10'd174) && (Y_Pos < 10'd217)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd190) && (X_Pos < 10'd194) && (Y_Pos > 10'd175) && (Y_Pos < 10'd217)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd449) && (Y_Pos > 10'd175) && (Y_Pos < 10'd217)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd279) && (X_Pos < 10'd283) && (Y_Pos > 10'd178) && (Y_Pos < 10'd183)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd313) && (X_Pos < 10'd317) && (Y_Pos > 10'd178) && (Y_Pos < 10'd183)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd322) && (X_Pos < 10'd326) && (Y_Pos > 10'd178) && (Y_Pos < 10'd183)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd356) && (X_Pos < 10'd360) && (Y_Pos > 10'd178) && (Y_Pos < 10'd183)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd278) && (X_Pos < 10'd282) && (Y_Pos > 10'd179) && (Y_Pos < 10'd184)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd314) && (X_Pos < 10'd318) && (Y_Pos > 10'd179) && (Y_Pos < 10'd184)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd321) && (X_Pos < 10'd325) && (Y_Pos > 10'd179) && (Y_Pos < 10'd184)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd357) && (X_Pos < 10'd361) && (Y_Pos > 10'd179) && (Y_Pos < 10'd184)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd241) && (X_Pos < 10'd281) && (Y_Pos > 10'd180) && (Y_Pos < 10'd185)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd315) && (X_Pos < 10'd324) && (Y_Pos > 10'd180) && (Y_Pos < 10'd185)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd358) && (X_Pos < 10'd398) && (Y_Pos > 10'd180) && (Y_Pos < 10'd185)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd240) && (X_Pos < 10'd244) && (Y_Pos > 10'd181) && (Y_Pos < 10'd186)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd395) && (X_Pos < 10'd399) && (Y_Pos > 10'd181) && (Y_Pos < 10'd186)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd239) && (X_Pos < 10'd243) && (Y_Pos > 10'd182) && (Y_Pos < 10'd219)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd400) && (Y_Pos > 10'd182) && (Y_Pos < 10'd219)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd242) && (Y_Pos > 10'd183) && (Y_Pos < 10'd220)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd397) && (X_Pos < 10'd401) && (Y_Pos > 10'd183) && (Y_Pos < 10'd220)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd237) && (X_Pos < 10'd241) && (Y_Pos > 10'd184) && (Y_Pos < 10'd188)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd398) && (X_Pos < 10'd402) && (Y_Pos > 10'd184) && (Y_Pos < 10'd188)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd270) && (X_Pos < 10'd305) && (Y_Pos > 10'd207) && (Y_Pos < 10'd212)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd334) && (X_Pos < 10'd369) && (Y_Pos > 10'd207) && (Y_Pos < 10'd212)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd302) && (X_Pos < 10'd306) && (Y_Pos > 10'd207) && (Y_Pos < 10'd217)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd333) && (X_Pos < 10'd337) && (Y_Pos > 10'd207) && (Y_Pos < 10'd217)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd207) && (Y_Pos < 10'd262)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd207) && (Y_Pos < 10'd262)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd303) && (X_Pos < 10'd307) && (Y_Pos > 10'd208) && (Y_Pos < 10'd216)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd332) && (X_Pos < 10'd336) && (Y_Pos > 10'd208) && (Y_Pos < 10'd216)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd304) && (X_Pos < 10'd335) && (Y_Pos > 10'd209) && (Y_Pos < 10'd215)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd275) && (X_Pos < 10'd305) && (Y_Pos > 10'd212) && (Y_Pos < 10'd217)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd334) && (X_Pos < 10'd364) && (Y_Pos > 10'd212) && (Y_Pos < 10'd217)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd274) && (X_Pos < 10'd278) && (Y_Pos > 10'd212) && (Y_Pos < 10'd257)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd361) && (X_Pos < 10'd365) && (Y_Pos > 10'd212) && (Y_Pos < 10'd257)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd273) && (X_Pos < 10'd277) && (Y_Pos > 10'd213) && (Y_Pos < 10'd257)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd362) && (X_Pos < 10'd366) && (Y_Pos > 10'd213) && (Y_Pos < 10'd257)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd185) && (X_Pos < 10'd190) && (Y_Pos > 10'd214) && (Y_Pos < 10'd218)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd449) && (X_Pos < 10'd454) && (Y_Pos > 10'd214) && (Y_Pos < 10'd218)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd188) && (Y_Pos > 10'd214) && (Y_Pos < 10'd219)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd187) && (X_Pos < 10'd192) && (Y_Pos > 10'd214) && (Y_Pos < 10'd219)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd447) && (X_Pos < 10'd452) && (Y_Pos > 10'd214) && (Y_Pos < 10'd219)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd451) && (X_Pos < 10'd521) && (Y_Pos > 10'd214) && (Y_Pos < 10'd219)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd237) && (X_Pos < 10'd241) && (Y_Pos > 10'd216) && (Y_Pos < 10'd221)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd398) && (X_Pos < 10'd402) && (Y_Pos > 10'd216) && (Y_Pos < 10'd221)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd194) && (X_Pos < 10'd198) && (Y_Pos > 10'd217) && (Y_Pos < 10'd221)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd441) && (X_Pos < 10'd445) && (Y_Pos > 10'd217) && (Y_Pos < 10'd221)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd193) && (X_Pos < 10'd197) && (Y_Pos > 10'd217) && (Y_Pos < 10'd222)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd227) && (X_Pos < 10'd232) && (Y_Pos > 10'd217) && (Y_Pos < 10'd222)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd236) && (X_Pos < 10'd240) && (Y_Pos > 10'd217) && (Y_Pos < 10'd222)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd399) && (X_Pos < 10'd403) && (Y_Pos > 10'd217) && (Y_Pos < 10'd222)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd407) && (X_Pos < 10'd412) && (Y_Pos > 10'd217) && (Y_Pos < 10'd222)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd442) && (X_Pos < 10'd446) && (Y_Pos > 10'd217) && (Y_Pos < 10'd222)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd196) && (Y_Pos > 10'd218) && (Y_Pos < 10'd223)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd229) && (X_Pos < 10'd239) && (Y_Pos > 10'd218) && (Y_Pos < 10'd223)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd400) && (X_Pos < 10'd410) && (Y_Pos > 10'd218) && (Y_Pos < 10'd223)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd443) && (X_Pos < 10'd521) && (Y_Pos > 10'd218) && (Y_Pos < 10'd223)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd196) && (Y_Pos > 10'd246) && (Y_Pos < 10'd251)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd229) && (X_Pos < 10'd239) && (Y_Pos > 10'd246) && (Y_Pos < 10'd251)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd400) && (X_Pos < 10'd410) && (Y_Pos > 10'd246) && (Y_Pos < 10'd251)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd443) && (X_Pos < 10'd521) && (Y_Pos > 10'd246) && (Y_Pos < 10'd251)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd193) && (X_Pos < 10'd197) && (Y_Pos > 10'd247) && (Y_Pos < 10'd252)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd228) && (X_Pos < 10'd232) && (Y_Pos > 10'd247) && (Y_Pos < 10'd252)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd236) && (X_Pos < 10'd240) && (Y_Pos > 10'd247) && (Y_Pos < 10'd252)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd399) && (X_Pos < 10'd403) && (Y_Pos > 10'd247) && (Y_Pos < 10'd252)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd407) && (X_Pos < 10'd411) && (Y_Pos > 10'd247) && (Y_Pos < 10'd252)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd442) && (X_Pos < 10'd446) && (Y_Pos > 10'd247) && (Y_Pos < 10'd252)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd227) && (X_Pos < 10'd231) && (Y_Pos > 10'd248) && (Y_Pos < 10'd252)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd408) && (X_Pos < 10'd412) && (Y_Pos > 10'd248) && (Y_Pos < 10'd252)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd194) && (X_Pos < 10'd198) && (Y_Pos > 10'd248) && (Y_Pos < 10'd253)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd237) && (X_Pos < 10'd241) && (Y_Pos > 10'd248) && (Y_Pos < 10'd253)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd398) && (X_Pos < 10'd402) && (Y_Pos > 10'd248) && (Y_Pos < 10'd253)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd441) && (X_Pos < 10'd445) && (Y_Pos > 10'd248) && (Y_Pos < 10'd253)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd199) && (Y_Pos > 10'd249) && (Y_Pos < 10'd297)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd229) && (Y_Pos > 10'd249) && (Y_Pos < 10'd297)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd242) && (Y_Pos > 10'd249) && (Y_Pos < 10'd297)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd397) && (X_Pos < 10'd401) && (Y_Pos > 10'd249) && (Y_Pos < 10'd297)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd410) && (X_Pos < 10'd414) && (Y_Pos > 10'd249) && (Y_Pos < 10'd297)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd440) && (X_Pos < 10'd444) && (Y_Pos > 10'd249) && (Y_Pos < 10'd297)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd226) && (X_Pos < 10'd230) && (Y_Pos > 10'd249) && (Y_Pos < 10'd298)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd413) && (Y_Pos > 10'd249) && (Y_Pos < 10'd298)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd196) && (X_Pos < 10'd200) && (Y_Pos > 10'd250) && (Y_Pos < 10'd297)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd239) && (X_Pos < 10'd243) && (Y_Pos > 10'd250) && (Y_Pos < 10'd297)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd400) && (Y_Pos > 10'd250) && (Y_Pos < 10'd297)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd443) && (Y_Pos > 10'd250) && (Y_Pos < 10'd297)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd192) && (Y_Pos > 10'd251) && (Y_Pos < 10'd256)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd447) && (X_Pos < 10'd521) && (Y_Pos > 10'd251) && (Y_Pos < 10'd256)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd275) && (X_Pos < 10'd364) && (Y_Pos > 10'd252) && (Y_Pos < 10'd257)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd190) && (X_Pos < 10'd194) && (Y_Pos > 10'd252) && (Y_Pos < 10'd294)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd445) && (X_Pos < 10'd449) && (Y_Pos > 10'd252) && (Y_Pos < 10'd294)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd189) && (X_Pos < 10'd193) && (Y_Pos > 10'd252) && (Y_Pos < 10'd295)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd446) && (X_Pos < 10'd450) && (Y_Pos > 10'd252) && (Y_Pos < 10'd295)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd270) && (X_Pos < 10'd369) && (Y_Pos > 10'd257) && (Y_Pos < 10'd262)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd272) && (X_Pos < 10'd367) && (Y_Pos > 10'd285) && (Y_Pos < 10'd289)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd270) && (X_Pos < 10'd275) && (Y_Pos > 10'd286) && (Y_Pos < 10'd291)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd364) && (X_Pos < 10'd369) && (Y_Pos > 10'd286) && (Y_Pos < 10'd291)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd272) && (Y_Pos > 10'd288) && (Y_Pos < 10'd297)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd367) && (X_Pos < 10'd371) && (Y_Pos > 10'd288) && (Y_Pos < 10'd297)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd269) && (X_Pos < 10'd273) && (Y_Pos > 10'd288) && (Y_Pos < 10'd298)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd370) && (Y_Pos > 10'd288) && (Y_Pos < 10'd298)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd125) && (X_Pos < 10'd192) && (Y_Pos > 10'd291) && (Y_Pos < 10'd296)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd447) && (X_Pos < 10'd514) && (Y_Pos > 10'd291) && (Y_Pos < 10'd296)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd124) && (X_Pos < 10'd128) && (Y_Pos > 10'd293) && (Y_Pos < 10'd297)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd515) && (Y_Pos > 10'd293) && (Y_Pos < 10'd297)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd122) && (X_Pos < 10'd127) && (Y_Pos > 10'd293) && (Y_Pos < 10'd298)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd512) && (X_Pos < 10'd517) && (Y_Pos > 10'd293) && (Y_Pos < 10'd298)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd193) && (X_Pos < 10'd198) && (Y_Pos > 10'd294) && (Y_Pos < 10'd299)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd227) && (X_Pos < 10'd231) && (Y_Pos > 10'd294) && (Y_Pos < 10'd299)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd236) && (X_Pos < 10'd241) && (Y_Pos > 10'd294) && (Y_Pos < 10'd299)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd270) && (X_Pos < 10'd274) && (Y_Pos > 10'd294) && (Y_Pos < 10'd299)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd365) && (X_Pos < 10'd369) && (Y_Pos > 10'd294) && (Y_Pos < 10'd299)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd398) && (X_Pos < 10'd403) && (Y_Pos > 10'd294) && (Y_Pos < 10'd299)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd408) && (X_Pos < 10'd412) && (Y_Pos > 10'd294) && (Y_Pos < 10'd299)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd441) && (X_Pos < 10'd446) && (Y_Pos > 10'd294) && (Y_Pos < 10'd299)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd121) && (X_Pos < 10'd125) && (Y_Pos > 10'd294) && (Y_Pos < 10'd300)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd514) && (X_Pos < 10'd518) && (Y_Pos > 10'd294) && (Y_Pos < 10'd300)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd120) && (X_Pos < 10'd124) && (Y_Pos > 10'd294) && (Y_Pos < 10'd301)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd515) && (X_Pos < 10'd519) && (Y_Pos > 10'd294) && (Y_Pos < 10'd301)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd228) && (X_Pos < 10'd232) && (Y_Pos > 10'd295) && (Y_Pos < 10'd299)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd407) && (X_Pos < 10'd411) && (Y_Pos > 10'd295) && (Y_Pos < 10'd299)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd271) && (X_Pos < 10'd275) && (Y_Pos > 10'd295) && (Y_Pos < 10'd300)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd364) && (X_Pos < 10'd368) && (Y_Pos > 10'd295) && (Y_Pos < 10'd300)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd235) && (X_Pos < 10'd239) && (Y_Pos > 10'd296) && (Y_Pos < 10'd300)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd400) && (X_Pos < 10'd404) && (Y_Pos > 10'd296) && (Y_Pos < 10'd300)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd127) && (X_Pos < 10'd196) && (Y_Pos > 10'd296) && (Y_Pos < 10'd301)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd229) && (X_Pos < 10'd238) && (Y_Pos > 10'd296) && (Y_Pos < 10'd301)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd272) && (X_Pos < 10'd312) && (Y_Pos > 10'd296) && (Y_Pos < 10'd301)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd327) && (X_Pos < 10'd367) && (Y_Pos > 10'd296) && (Y_Pos < 10'd301)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd401) && (X_Pos < 10'd410) && (Y_Pos > 10'd296) && (Y_Pos < 10'd301)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd443) && (X_Pos < 10'd512) && (Y_Pos > 10'd296) && (Y_Pos < 10'd301)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd126) && (X_Pos < 10'd130) && (Y_Pos > 10'd297) && (Y_Pos < 10'd302)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd309) && (X_Pos < 10'd313) && (Y_Pos > 10'd297) && (Y_Pos < 10'd302)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd326) && (X_Pos < 10'd330) && (Y_Pos > 10'd297) && (Y_Pos < 10'd302)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd509) && (X_Pos < 10'd513) && (Y_Pos > 10'd297) && (Y_Pos < 10'd302)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd125) && (X_Pos < 10'd129) && (Y_Pos > 10'd298) && (Y_Pos < 10'd303)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd310) && (X_Pos < 10'd314) && (Y_Pos > 10'd298) && (Y_Pos < 10'd303)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd325) && (X_Pos < 10'd329) && (Y_Pos > 10'd298) && (Y_Pos < 10'd303)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd510) && (X_Pos < 10'd514) && (Y_Pos > 10'd298) && (Y_Pos < 10'd303)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd118) && (X_Pos < 10'd123) && (Y_Pos > 10'd298) && (Y_Pos < 10'd443)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd516) && (X_Pos < 10'd521) && (Y_Pos > 10'd298) && (Y_Pos < 10'd443)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd315) && (Y_Pos > 10'd299) && (Y_Pos < 10'd336)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd324) && (X_Pos < 10'd328) && (Y_Pos > 10'd299) && (Y_Pos < 10'd336)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd127) && (Y_Pos > 10'd299) && (Y_Pos < 10'd363)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd512) && (X_Pos < 10'd516) && (Y_Pos > 10'd299) && (Y_Pos < 10'd363)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd124) && (X_Pos < 10'd128) && (Y_Pos > 10'd299) && (Y_Pos < 10'd364)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd515) && (Y_Pos > 10'd299) && (Y_Pos < 10'd364)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd312) && (X_Pos < 10'd316) && (Y_Pos > 10'd300) && (Y_Pos < 10'd337)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd327) && (Y_Pos > 10'd300) && (Y_Pos < 10'd337)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd158) && (X_Pos < 10'd196) && (Y_Pos > 10'd323) && (Y_Pos < 10'd328)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd229) && (X_Pos < 10'd281) && (Y_Pos > 10'd323) && (Y_Pos < 10'd328)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd358) && (X_Pos < 10'd410) && (Y_Pos > 10'd323) && (Y_Pos < 10'd328)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd443) && (X_Pos < 10'd481) && (Y_Pos > 10'd323) && (Y_Pos < 10'd328)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd157) && (X_Pos < 10'd161) && (Y_Pos > 10'd324) && (Y_Pos < 10'd329)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd278) && (X_Pos < 10'd282) && (Y_Pos > 10'd324) && (Y_Pos < 10'd329)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd357) && (X_Pos < 10'd361) && (Y_Pos > 10'd324) && (Y_Pos < 10'd329)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd478) && (X_Pos < 10'd482) && (Y_Pos > 10'd324) && (Y_Pos < 10'd329)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd228) && (X_Pos < 10'd232) && (Y_Pos > 10'd325) && (Y_Pos < 10'd329)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd407) && (X_Pos < 10'd411) && (Y_Pos > 10'd325) && (Y_Pos < 10'd329)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd156) && (X_Pos < 10'd160) && (Y_Pos > 10'd325) && (Y_Pos < 10'd330)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd193) && (X_Pos < 10'd198) && (Y_Pos > 10'd325) && (Y_Pos < 10'd330)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd227) && (X_Pos < 10'd231) && (Y_Pos > 10'd325) && (Y_Pos < 10'd330)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd279) && (X_Pos < 10'd283) && (Y_Pos > 10'd325) && (Y_Pos < 10'd330)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd356) && (X_Pos < 10'd360) && (Y_Pos > 10'd325) && (Y_Pos < 10'd330)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd408) && (X_Pos < 10'd412) && (Y_Pos > 10'd325) && (Y_Pos < 10'd330)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd441) && (X_Pos < 10'd446) && (Y_Pos > 10'd325) && (Y_Pos < 10'd330)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd479) && (X_Pos < 10'd483) && (Y_Pos > 10'd325) && (Y_Pos < 10'd330)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd226) && (X_Pos < 10'd230) && (Y_Pos > 10'd326) && (Y_Pos < 10'd336)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd413) && (Y_Pos > 10'd326) && (Y_Pos < 10'd336)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd155) && (X_Pos < 10'd159) && (Y_Pos > 10'd326) && (Y_Pos < 10'd337)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd280) && (X_Pos < 10'd284) && (Y_Pos > 10'd326) && (Y_Pos < 10'd337)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd355) && (X_Pos < 10'd359) && (Y_Pos > 10'd326) && (Y_Pos < 10'd337)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd480) && (X_Pos < 10'd484) && (Y_Pos > 10'd326) && (Y_Pos < 10'd337)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd154) && (X_Pos < 10'd158) && (Y_Pos > 10'd327) && (Y_Pos < 10'd336)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd229) && (Y_Pos > 10'd327) && (Y_Pos < 10'd336)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd281) && (X_Pos < 10'd285) && (Y_Pos > 10'd327) && (Y_Pos < 10'd336)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd354) && (X_Pos < 10'd358) && (Y_Pos > 10'd327) && (Y_Pos < 10'd336)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd410) && (X_Pos < 10'd414) && (Y_Pos > 10'd327) && (Y_Pos < 10'd336)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd481) && (X_Pos < 10'd485) && (Y_Pos > 10'd327) && (Y_Pos < 10'd336)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd196) && (X_Pos < 10'd200) && (Y_Pos > 10'd327) && (Y_Pos < 10'd374)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd439) && (X_Pos < 10'd443) && (Y_Pos > 10'd327) && (Y_Pos < 10'd374)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd195) && (X_Pos < 10'd199) && (Y_Pos > 10'd327) && (Y_Pos < 10'd375)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd440) && (X_Pos < 10'd444) && (Y_Pos > 10'd327) && (Y_Pos < 10'd375)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd156) && (X_Pos < 10'd160) && (Y_Pos > 10'd333) && (Y_Pos < 10'd338)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd227) && (X_Pos < 10'd232) && (Y_Pos > 10'd333) && (Y_Pos < 10'd338)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd279) && (X_Pos < 10'd283) && (Y_Pos > 10'd333) && (Y_Pos < 10'd338)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd313) && (X_Pos < 10'd317) && (Y_Pos > 10'd333) && (Y_Pos < 10'd338)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd322) && (X_Pos < 10'd326) && (Y_Pos > 10'd333) && (Y_Pos < 10'd338)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd356) && (X_Pos < 10'd360) && (Y_Pos > 10'd333) && (Y_Pos < 10'd338)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd407) && (X_Pos < 10'd412) && (Y_Pos > 10'd333) && (Y_Pos < 10'd338)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd479) && (X_Pos < 10'd483) && (Y_Pos > 10'd333) && (Y_Pos < 10'd338)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd157) && (X_Pos < 10'd161) && (Y_Pos > 10'd334) && (Y_Pos < 10'd339)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd278) && (X_Pos < 10'd282) && (Y_Pos > 10'd334) && (Y_Pos < 10'd339)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd314) && (X_Pos < 10'd318) && (Y_Pos > 10'd334) && (Y_Pos < 10'd339)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd321) && (X_Pos < 10'd325) && (Y_Pos > 10'd334) && (Y_Pos < 10'd339)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd357) && (X_Pos < 10'd361) && (Y_Pos > 10'd334) && (Y_Pos < 10'd339)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd478) && (X_Pos < 10'd482) && (Y_Pos > 10'd334) && (Y_Pos < 10'd339)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd158) && (X_Pos < 10'd183) && (Y_Pos > 10'd335) && (Y_Pos < 10'd339)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd229) && (X_Pos < 10'd281) && (Y_Pos > 10'd335) && (Y_Pos < 10'd339)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd315) && (X_Pos < 10'd324) && (Y_Pos > 10'd335) && (Y_Pos < 10'd339)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd358) && (X_Pos < 10'd410) && (Y_Pos > 10'd335) && (Y_Pos < 10'd339)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd456) && (X_Pos < 10'd481) && (Y_Pos > 10'd335) && (Y_Pos < 10'd339)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd180) && (X_Pos < 10'd184) && (Y_Pos > 10'd336) && (Y_Pos < 10'd340)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd455) && (X_Pos < 10'd459) && (Y_Pos > 10'd336) && (Y_Pos < 10'd340)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd181) && (X_Pos < 10'd185) && (Y_Pos > 10'd336) && (Y_Pos < 10'd341)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd454) && (X_Pos < 10'd458) && (Y_Pos > 10'd336) && (Y_Pos < 10'd341)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd182) && (X_Pos < 10'd186) && (Y_Pos > 10'd337) && (Y_Pos < 10'd375)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd453) && (X_Pos < 10'd457) && (Y_Pos > 10'd337) && (Y_Pos < 10'd375)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd183) && (X_Pos < 10'd187) && (Y_Pos > 10'd338) && (Y_Pos < 10'd375)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd452) && (X_Pos < 10'd456) && (Y_Pos > 10'd338) && (Y_Pos < 10'd375)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd125) && (X_Pos < 10'd129) && (Y_Pos > 10'd360) && (Y_Pos < 10'd365)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd510) && (X_Pos < 10'd514) && (Y_Pos > 10'd360) && (Y_Pos < 10'd365)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd126) && (X_Pos < 10'd130) && (Y_Pos > 10'd361) && (Y_Pos < 10'd365)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd509) && (X_Pos < 10'd513) && (Y_Pos > 10'd361) && (Y_Pos < 10'd365)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd127) && (X_Pos < 10'd153) && (Y_Pos > 10'd362) && (Y_Pos < 10'd367)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd229) && (X_Pos < 10'd239) && (Y_Pos > 10'd362) && (Y_Pos < 10'd367)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd272) && (X_Pos < 10'd367) && (Y_Pos > 10'd362) && (Y_Pos < 10'd367)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd400) && (X_Pos < 10'd410) && (Y_Pos > 10'd362) && (Y_Pos < 10'd367)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd486) && (X_Pos < 10'd512) && (Y_Pos > 10'd362) && (Y_Pos < 10'd367)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd150) && (X_Pos < 10'd154) && (Y_Pos > 10'd363) && (Y_Pos < 10'd368)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd228) && (X_Pos < 10'd232) && (Y_Pos > 10'd363) && (Y_Pos < 10'd368)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd271) && (X_Pos < 10'd275) && (Y_Pos > 10'd363) && (Y_Pos < 10'd368)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd364) && (X_Pos < 10'd368) && (Y_Pos > 10'd363) && (Y_Pos < 10'd368)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd407) && (X_Pos < 10'd411) && (Y_Pos > 10'd363) && (Y_Pos < 10'd368)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd485) && (X_Pos < 10'd489) && (Y_Pos > 10'd363) && (Y_Pos < 10'd368)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd236) && (X_Pos < 10'd240) && (Y_Pos > 10'd364) && (Y_Pos < 10'd368)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd399) && (X_Pos < 10'd403) && (Y_Pos > 10'd364) && (Y_Pos < 10'd368)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd151) && (X_Pos < 10'd155) && (Y_Pos > 10'd364) && (Y_Pos < 10'd369)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd227) && (X_Pos < 10'd231) && (Y_Pos > 10'd364) && (Y_Pos < 10'd369)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd237) && (X_Pos < 10'd241) && (Y_Pos > 10'd364) && (Y_Pos < 10'd369)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd270) && (X_Pos < 10'd274) && (Y_Pos > 10'd364) && (Y_Pos < 10'd369)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd365) && (X_Pos < 10'd369) && (Y_Pos > 10'd364) && (Y_Pos < 10'd369)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd398) && (X_Pos < 10'd402) && (Y_Pos > 10'd364) && (Y_Pos < 10'd369)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd408) && (X_Pos < 10'd412) && (Y_Pos > 10'd364) && (Y_Pos < 10'd369)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd484) && (X_Pos < 10'd488) && (Y_Pos > 10'd364) && (Y_Pos < 10'd369)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd152) && (X_Pos < 10'd156) && (Y_Pos > 10'd365) && (Y_Pos < 10'd375)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd268) && (X_Pos < 10'd273) && (Y_Pos > 10'd365) && (Y_Pos < 10'd375)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd366) && (X_Pos < 10'd371) && (Y_Pos > 10'd365) && (Y_Pos < 10'd375)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd483) && (X_Pos < 10'd487) && (Y_Pos > 10'd365) && (Y_Pos < 10'd375)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd226) && (X_Pos < 10'd230) && (Y_Pos > 10'd365) && (Y_Pos < 10'd402)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd238) && (X_Pos < 10'd242) && (Y_Pos > 10'd365) && (Y_Pos < 10'd402)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd397) && (X_Pos < 10'd401) && (Y_Pos > 10'd365) && (Y_Pos < 10'd402)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd409) && (X_Pos < 10'd413) && (Y_Pos > 10'd365) && (Y_Pos < 10'd402)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd225) && (X_Pos < 10'd229) && (Y_Pos > 10'd365) && (Y_Pos < 10'd403)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd410) && (X_Pos < 10'd414) && (Y_Pos > 10'd365) && (Y_Pos < 10'd403)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd153) && (X_Pos < 10'd157) && (Y_Pos > 10'd366) && (Y_Pos < 10'd375)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd482) && (X_Pos < 10'd486) && (Y_Pos > 10'd366) && (Y_Pos < 10'd375)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd239) && (X_Pos < 10'd243) && (Y_Pos > 10'd366) && (Y_Pos < 10'd403)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd396) && (X_Pos < 10'd400) && (Y_Pos > 10'd366) && (Y_Pos < 10'd403)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd151) && (X_Pos < 10'd155) && (Y_Pos > 10'd371) && (Y_Pos < 10'd376)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd184) && (X_Pos < 10'd188) && (Y_Pos > 10'd371) && (Y_Pos < 10'd376)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd194) && (X_Pos < 10'd198) && (Y_Pos > 10'd371) && (Y_Pos < 10'd376)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd441) && (X_Pos < 10'd445) && (Y_Pos > 10'd371) && (Y_Pos < 10'd376)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd451) && (X_Pos < 10'd455) && (Y_Pos > 10'd371) && (Y_Pos < 10'd376)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd484) && (X_Pos < 10'd488) && (Y_Pos > 10'd371) && (Y_Pos < 10'd376)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd150) && (X_Pos < 10'd154) && (Y_Pos > 10'd372) && (Y_Pos < 10'd377)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd185) && (X_Pos < 10'd189) && (Y_Pos > 10'd372) && (Y_Pos < 10'd377)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd193) && (X_Pos < 10'd197) && (Y_Pos > 10'd372) && (Y_Pos < 10'd377)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd270) && (X_Pos < 10'd275) && (Y_Pos > 10'd372) && (Y_Pos < 10'd377)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd364) && (X_Pos < 10'd369) && (Y_Pos > 10'd372) && (Y_Pos < 10'd377)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd442) && (X_Pos < 10'd446) && (Y_Pos > 10'd372) && (Y_Pos < 10'd377)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd450) && (X_Pos < 10'd454) && (Y_Pos > 10'd372) && (Y_Pos < 10'd377)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd485) && (X_Pos < 10'd489) && (Y_Pos > 10'd372) && (Y_Pos < 10'd377)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd127) && (X_Pos < 10'd153) && (Y_Pos > 10'd373) && (Y_Pos < 10'd378)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd186) && (X_Pos < 10'd196) && (Y_Pos > 10'd373) && (Y_Pos < 10'd378)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd272) && (X_Pos < 10'd312) && (Y_Pos > 10'd373) && (Y_Pos < 10'd378)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd327) && (X_Pos < 10'd367) && (Y_Pos > 10'd373) && (Y_Pos < 10'd378)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd443) && (X_Pos < 10'd453) && (Y_Pos > 10'd373) && (Y_Pos < 10'd378)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd486) && (X_Pos < 10'd512) && (Y_Pos > 10'd373) && (Y_Pos < 10'd378)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd125) && (X_Pos < 10'd130) && (Y_Pos > 10'd375) && (Y_Pos < 10'd380)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd309) && (X_Pos < 10'd314) && (Y_Pos > 10'd375) && (Y_Pos < 10'd380)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd325) && (X_Pos < 10'd330) && (Y_Pos > 10'd375) && (Y_Pos < 10'd380)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd509) && (X_Pos < 10'd514) && (Y_Pos > 10'd375) && (Y_Pos < 10'd380)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd311) && (X_Pos < 10'd315) && (Y_Pos > 10'd377) && (Y_Pos < 10'd413)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd324) && (X_Pos < 10'd328) && (Y_Pos > 10'd377) && (Y_Pos < 10'd413)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd312) && (X_Pos < 10'd316) && (Y_Pos > 10'd377) && (Y_Pos < 10'd414)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd323) && (X_Pos < 10'd327) && (Y_Pos > 10'd377) && (Y_Pos < 10'd414)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd123) && (X_Pos < 10'd128) && (Y_Pos > 10'd377) && (Y_Pos < 10'd441)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd516) && (Y_Pos > 10'd377) && (Y_Pos < 10'd441)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd237) && (X_Pos < 10'd241) && (Y_Pos > 10'd397) && (Y_Pos < 10'd401)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd398) && (X_Pos < 10'd402) && (Y_Pos > 10'd397) && (Y_Pos < 10'd401)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd223) && (X_Pos < 10'd228) && (Y_Pos > 10'd399) && (Y_Pos < 10'd404)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd240) && (X_Pos < 10'd244) && (Y_Pos > 10'd399) && (Y_Pos < 10'd404)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd395) && (X_Pos < 10'd399) && (Y_Pos > 10'd399) && (Y_Pos < 10'd404)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd411) && (X_Pos < 10'd416) && (Y_Pos > 10'd399) && (Y_Pos < 10'd404)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd241) && (X_Pos < 10'd245) && (Y_Pos > 10'd400) && (Y_Pos < 10'd405)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd394) && (X_Pos < 10'd398) && (Y_Pos > 10'd400) && (Y_Pos < 10'd405)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd157) && (X_Pos < 10'd226) && (Y_Pos > 10'd401) && (Y_Pos < 10'd406)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd242) && (X_Pos < 10'd282) && (Y_Pos > 10'd401) && (Y_Pos < 10'd406)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd357) && (X_Pos < 10'd397) && (Y_Pos > 10'd401) && (Y_Pos < 10'd406)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd413) && (X_Pos < 10'd482) && (Y_Pos > 10'd401) && (Y_Pos < 10'd406)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd156) && (X_Pos < 10'd160) && (Y_Pos > 10'd402) && (Y_Pos < 10'd407)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd279) && (X_Pos < 10'd283) && (Y_Pos > 10'd402) && (Y_Pos < 10'd407)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd356) && (X_Pos < 10'd360) && (Y_Pos > 10'd402) && (Y_Pos < 10'd407)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd479) && (X_Pos < 10'd483) && (Y_Pos > 10'd402) && (Y_Pos < 10'd407)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd155) && (X_Pos < 10'd159) && (Y_Pos > 10'd403) && (Y_Pos < 10'd415)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd280) && (X_Pos < 10'd284) && (Y_Pos > 10'd403) && (Y_Pos < 10'd415)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd355) && (X_Pos < 10'd359) && (Y_Pos > 10'd403) && (Y_Pos < 10'd415)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd480) && (X_Pos < 10'd484) && (Y_Pos > 10'd403) && (Y_Pos < 10'd415)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd154) && (X_Pos < 10'd158) && (Y_Pos > 10'd404) && (Y_Pos < 10'd413)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd281) && (X_Pos < 10'd285) && (Y_Pos > 10'd404) && (Y_Pos < 10'd413)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd354) && (X_Pos < 10'd358) && (Y_Pos > 10'd404) && (Y_Pos < 10'd413)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd481) && (X_Pos < 10'd485) && (Y_Pos > 10'd404) && (Y_Pos < 10'd413)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd156) && (X_Pos < 10'd160) && (Y_Pos > 10'd410) && (Y_Pos < 10'd415)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd279) && (X_Pos < 10'd283) && (Y_Pos > 10'd410) && (Y_Pos < 10'd415)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd313) && (X_Pos < 10'd317) && (Y_Pos > 10'd410) && (Y_Pos < 10'd415)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd322) && (X_Pos < 10'd326) && (Y_Pos > 10'd410) && (Y_Pos < 10'd415)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd356) && (X_Pos < 10'd360) && (Y_Pos > 10'd410) && (Y_Pos < 10'd415)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd479) && (X_Pos < 10'd483) && (Y_Pos > 10'd410) && (Y_Pos < 10'd415)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd314) && (X_Pos < 10'd318) && (Y_Pos > 10'd411) && (Y_Pos < 10'd416)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd321) && (X_Pos < 10'd325) && (Y_Pos > 10'd411) && (Y_Pos < 10'd416)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd157) && (X_Pos < 10'd161) && (Y_Pos > 10'd412) && (Y_Pos < 10'd416)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd278) && (X_Pos < 10'd282) && (Y_Pos > 10'd412) && (Y_Pos < 10'd416)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd357) && (X_Pos < 10'd361) && (Y_Pos > 10'd412) && (Y_Pos < 10'd416)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd478) && (X_Pos < 10'd482) && (Y_Pos > 10'd412) && (Y_Pos < 10'd416)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd158) && (X_Pos < 10'd281) && (Y_Pos > 10'd412) && (Y_Pos < 10'd417)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd315) && (X_Pos < 10'd324) && (Y_Pos > 10'd412) && (Y_Pos < 10'd417)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd358) && (X_Pos < 10'd481) && (Y_Pos > 10'd412) && (Y_Pos < 10'd417)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd125) && (X_Pos < 10'd130) && (Y_Pos > 10'd438) && (Y_Pos < 10'd443)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd509) && (X_Pos < 10'd514) && (Y_Pos > 10'd438) && (Y_Pos < 10'd443)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd127) && (X_Pos < 10'd512) && (Y_Pos > 10'd439) && (Y_Pos < 10'd444)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd120) && (X_Pos < 10'd125) && (Y_Pos > 10'd440) && (Y_Pos < 10'd446)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd514) && (X_Pos < 10'd519) && (Y_Pos > 10'd440) && (Y_Pos < 10'd446)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd122) && (X_Pos < 10'd128) && (Y_Pos > 10'd443) && (Y_Pos < 10'd447)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd511) && (X_Pos < 10'd517) && (Y_Pos > 10'd443) && (Y_Pos < 10'd447)) Is_Wall = 1'b1;

	if ((X_Pos > 10'd125) && (X_Pos < 10'd514) && (Y_Pos > 10'd444) && (Y_Pos < 10'd449)) Is_Wall = 1'b1;

	if (~Is_Wall) Is_Wall = 1'b0;
end

endmodule

